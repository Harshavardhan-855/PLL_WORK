* NGSPICE file created from vco.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_VC56GX a_1215_n800# a_63_n800# a_n1089_n800# a_n225_n800#
+ a_n1425_n897# a_399_831# a_1311_n800# a_927_n800# a_111_n897# a_n1185_n800# a_1263_n897#
+ a_879_n897# a_1359_831# a_n321_n800# a_n273_n897# a_15_831# a_n753_831# a_1023_n800#
+ a_639_n800# a_n1281_n800# a_591_831# a_n1233_n897# a_207_831# a_735_n800# a_n33_n800#
+ a_1071_n897# a_687_n897# a_n1469_n800# a_n897_n800# a_n945_831# a_831_n800# a_447_n800#
+ a_n81_n897# a_n849_n897# a_783_831# a_n993_n800# a_n1041_n897# a_543_n800# a_n177_831#
+ a_159_n800# a_n609_n800# a_495_n897# a_n1137_831# a_255_n800# a_n705_n800# a_975_831#
+ a_n657_n897# a_1407_n800# w_n1607_n1019# a_n369_831# a_351_n800# a_n417_n800# a_n801_n800#
+ a_n1329_831# a_1119_n800# a_n1377_n800# a_303_n897# a_1167_831# a_n129_n800# a_n513_n800#
+ a_n465_n897# a_n561_831#
X0 a_1023_n800# a_975_831# a_927_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1 a_n993_n800# a_n1041_n897# a_n1089_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2 a_n33_n800# a_n81_n897# a_n129_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3 a_351_n800# a_303_n897# a_255_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4 a_1311_n800# a_1263_n897# a_1215_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5 a_n1281_n800# a_n1329_831# a_n1377_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6 a_n609_n800# a_n657_n897# a_n705_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7 a_927_n800# a_879_n897# a_831_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8 a_n897_n800# a_n945_831# a_n993_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X9 a_255_n800# a_207_831# a_159_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X10 a_1215_n800# a_1167_831# a_1119_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X11 a_n321_n800# a_n369_831# a_n417_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X12 a_n1185_n800# a_n1233_n897# a_n1281_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X13 a_543_n800# a_495_n897# a_447_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X14 a_831_n800# a_783_831# a_735_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X15 a_159_n800# a_111_n897# a_63_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X16 a_1119_n800# a_1071_n897# a_1023_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X17 a_n225_n800# a_n273_n897# a_n321_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X18 a_n1089_n800# a_n1137_831# a_n1185_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X19 a_447_n800# a_399_831# a_351_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X20 a_1407_n800# a_1359_831# a_1311_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X21 a_n513_n800# a_n561_831# a_n609_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X22 a_63_n800# a_15_831# a_n33_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X23 a_735_n800# a_687_n897# a_639_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X24 a_n1377_n800# a_n1425_n897# a_n1469_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X25 a_n801_n800# a_n849_n897# a_n897_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X26 a_n129_n800# a_n177_831# a_n225_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X27 a_n417_n800# a_n465_n897# a_n513_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X28 a_639_n800# a_591_831# a_543_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X29 a_n705_n800# a_n753_831# a_n801_n800# w_n1607_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_UBPJLS a_n369_322# a_735_n300# a_n33_n300# a_n1329_322#
+ a_303_n388# a_n1469_n300# a_1167_322# a_n897_n300# a_n465_n388# a_n561_322# a_831_n300#
+ a_447_n300# a_n993_n300# a_n1425_n388# a_399_322# a_543_n300# a_159_n300# a_n609_n300#
+ a_879_n388# a_111_n388# a_1263_n388# a_1359_322# a_n753_322# a_15_322# a_n273_n388#
+ a_255_n300# a_n705_n300# a_1407_n300# a_591_322# a_n1233_n388# a_n1571_n474# a_351_n300#
+ a_n801_n300# a_207_322# a_n417_n300# a_1071_n388# a_687_n388# a_1119_n300# a_n1377_n300#
+ a_n945_322# a_n513_n300# a_n129_n300# a_783_322# a_n81_n388# a_n849_n388# a_1215_n300#
+ a_63_n300# a_n1089_n300# a_n177_322# a_n1041_n388# a_n225_n300# a_495_n388# a_1311_n300#
+ a_927_n300# a_n1185_n300# a_n1137_322# a_n321_n300# a_975_322# a_n657_n388# a_1023_n300#
+ a_639_n300# a_n1281_n300#
X0 a_n897_n300# a_n945_322# a_n993_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1 a_927_n300# a_879_n388# a_831_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X2 a_1215_n300# a_1167_322# a_1119_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X3 a_255_n300# a_207_322# a_159_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X4 a_n321_n300# a_n369_322# a_n417_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X5 a_543_n300# a_495_n388# a_447_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X6 a_n1185_n300# a_n1233_n388# a_n1281_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X7 a_831_n300# a_783_322# a_735_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X8 a_1119_n300# a_1071_n388# a_1023_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X9 a_159_n300# a_111_n388# a_63_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X10 a_n225_n300# a_n273_n388# a_n321_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X11 a_447_n300# a_399_322# a_351_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X12 a_1407_n300# a_1359_322# a_1311_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X13 a_n1089_n300# a_n1137_322# a_n1185_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X14 a_n513_n300# a_n561_322# a_n609_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X15 a_63_n300# a_15_322# a_n33_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X16 a_n1377_n300# a_n1425_n388# a_n1469_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X17 a_735_n300# a_687_n388# a_639_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X18 a_n801_n300# a_n849_n388# a_n897_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X19 a_n129_n300# a_n177_322# a_n225_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X20 a_n417_n300# a_n465_n388# a_n513_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X21 a_639_n300# a_591_322# a_543_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X22 a_n705_n300# a_n753_322# a_n801_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X23 a_1023_n300# a_975_322# a_927_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X24 a_1311_n300# a_1263_n388# a_1215_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X25 a_n993_n300# a_n1041_n388# a_n1089_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X26 a_n33_n300# a_n81_n388# a_n129_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X27 a_351_n300# a_303_n388# a_255_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X28 a_n1281_n300# a_n1329_322# a_n1377_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X29 a_n609_n300# a_n657_n388# a_n705_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_CDSMYA a_n369_322# a_735_n300# a_n33_n300# a_n1329_322#
+ a_303_n388# a_n1469_n300# a_1167_322# a_n897_n300# a_n465_n388# a_n561_322# a_831_n300#
+ a_447_n300# a_n993_n300# a_n1425_n388# a_399_322# a_543_n300# a_159_n300# a_n609_n300#
+ a_879_n388# a_111_n388# a_1263_n388# a_1359_322# a_n753_322# a_15_322# a_n273_n388#
+ a_255_n300# a_n705_n300# a_1407_n300# a_591_322# a_n1233_n388# a_n1571_n474# a_351_n300#
+ a_n801_n300# a_207_322# a_n417_n300# a_1071_n388# a_687_n388# a_1119_n300# a_n1377_n300#
+ a_n945_322# a_n513_n300# a_n129_n300# a_783_322# a_n81_n388# a_n849_n388# a_1215_n300#
+ a_63_n300# a_n1089_n300# a_n177_322# a_n1041_n388# a_n225_n300# a_495_n388# a_1311_n300#
+ a_927_n300# a_n1185_n300# a_n1137_322# a_n321_n300# a_975_322# a_n657_n388# a_1023_n300#
+ a_639_n300# a_n1281_n300#
X0 a_n897_n300# a_n945_322# a_n993_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1 a_927_n300# a_879_n388# a_831_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X2 a_1215_n300# a_1167_322# a_1119_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X3 a_255_n300# a_207_322# a_159_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X4 a_n321_n300# a_n369_322# a_n417_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X5 a_543_n300# a_495_n388# a_447_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X6 a_n1185_n300# a_n1233_n388# a_n1281_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X7 a_831_n300# a_783_322# a_735_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X8 a_1119_n300# a_1071_n388# a_1023_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X9 a_159_n300# a_111_n388# a_63_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X10 a_n225_n300# a_n273_n388# a_n321_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X11 a_447_n300# a_399_322# a_351_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X12 a_1407_n300# a_1359_322# a_1311_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X13 a_n1089_n300# a_n1137_322# a_n1185_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X14 a_n513_n300# a_n561_322# a_n609_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X15 a_63_n300# a_15_322# a_n33_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X16 a_n1377_n300# a_n1425_n388# a_n1469_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X17 a_735_n300# a_687_n388# a_639_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X18 a_n801_n300# a_n849_n388# a_n897_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X19 a_n129_n300# a_n177_322# a_n225_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X20 a_n417_n300# a_n465_n388# a_n513_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X21 a_639_n300# a_591_322# a_543_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X22 a_n705_n300# a_n753_322# a_n801_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X23 a_1023_n300# a_975_322# a_927_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X24 a_1311_n300# a_1263_n388# a_1215_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X25 a_n993_n300# a_n1041_n388# a_n1089_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X26 a_n33_n300# a_n81_n388# a_n129_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X27 a_351_n300# a_303_n388# a_255_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X28 a_n1281_n300# a_n1329_322# a_n1377_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X29 a_n609_n300# a_n657_n388# a_n705_n300# a_n1571_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_42S873 a_n81_n600# a_n269_n600# a_n129_622# a_n225_n688#
+ a_207_n600# a_n371_n774# a_n33_n688# a_15_n600# a_n177_n600# a_111_n600# a_159_n688#
+ a_63_622#
X0 a_n177_n600# a_n225_n688# a_n269_n600# a_n371_n774# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=1.86 ps=12.62 w=6 l=0.15
X1 a_207_n600# a_159_n688# a_111_n600# a_n371_n774# sky130_fd_pr__nfet_01v8 ad=1.86 pd=12.62 as=0.99 ps=6.33 w=6 l=0.15
X2 a_111_n600# a_63_622# a_15_n600# a_n371_n774# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.15
X3 a_n81_n600# a_n129_622# a_n177_n600# a_n371_n774# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.15
X4 a_15_n600# a_n33_n688# a_n81_n600# a_n371_n774# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_UYM7GH a_207_n1800# a_111_n1800# a_n81_n1800# a_n177_n1800#
+ a_n33_n1897# w_n407_n2019# a_n225_n1897# a_159_n1897# a_15_n1800# a_n129_1831# a_n269_n1800#
+ a_63_1831#
X0 a_n81_n1800# a_n129_1831# a_n177_n1800# w_n407_n2019# sky130_fd_pr__pfet_01v8 ad=2.97 pd=18.33 as=2.97 ps=18.33 w=18 l=0.15
X1 a_15_n1800# a_n33_n1897# a_n81_n1800# w_n407_n2019# sky130_fd_pr__pfet_01v8 ad=2.97 pd=18.33 as=2.97 ps=18.33 w=18 l=0.15
X2 a_n177_n1800# a_n225_n1897# a_n269_n1800# w_n407_n2019# sky130_fd_pr__pfet_01v8 ad=2.97 pd=18.33 as=5.58 ps=36.62 w=18 l=0.15
X3 a_111_n1800# a_63_1831# a_15_n1800# w_n407_n2019# sky130_fd_pr__pfet_01v8 ad=2.97 pd=18.33 as=2.97 ps=18.33 w=18 l=0.15
X4 a_207_n1800# a_159_n1897# a_111_n1800# w_n407_n2019# sky130_fd_pr__pfet_01v8 ad=5.58 pd=36.62 as=2.97 ps=18.33 w=18 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_VC5S4W w_n647_n1019# a_63_n800# a_n225_n800# a_399_831#
+ a_111_n897# a_n321_n800# a_n273_n897# a_15_831# a_207_831# a_n33_n800# a_n509_n800#
+ a_447_n800# a_n81_n897# a_n177_831# a_159_n800# a_255_n800# a_n369_831# a_351_n800#
+ a_n417_n800# a_303_n897# a_n129_n800# a_n465_n897#
X0 a_n33_n800# a_n81_n897# a_n129_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1 a_351_n800# a_303_n897# a_255_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2 a_255_n800# a_207_831# a_159_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3 a_n321_n800# a_n369_831# a_n417_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4 a_159_n800# a_111_n897# a_63_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5 a_n225_n800# a_n273_n897# a_n321_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6 a_447_n800# a_399_831# a_351_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X7 a_63_n800# a_15_831# a_n33_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8 a_n129_n800# a_n177_831# a_n225_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X9 a_n417_n800# a_n465_n897# a_n509_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_JT8PYA a_n369_322# a_n33_n300# a_n509_n300# a_303_n388#
+ a_n465_n388# a_447_n300# a_399_322# a_159_n300# a_111_n388# a_15_322# a_n273_n388#
+ a_255_n300# a_n611_n474# a_351_n300# a_207_322# a_n417_n300# a_n129_n300# a_n81_n388#
+ a_63_n300# a_n177_322# a_n225_n300# a_n321_n300#
X0 a_255_n300# a_207_322# a_159_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1 a_n321_n300# a_n369_322# a_n417_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X2 a_159_n300# a_111_n388# a_63_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X3 a_n225_n300# a_n273_n388# a_n321_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X4 a_447_n300# a_399_322# a_351_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X5 a_63_n300# a_15_322# a_n33_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X6 a_n129_n300# a_n177_322# a_n225_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X7 a_n417_n300# a_n465_n388# a_n509_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X8 a_n33_n300# a_n81_n388# a_n129_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X9 a_351_n300# a_303_n388# a_255_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_JLF2PR a_n369_322# a_n33_n300# a_n509_n300# a_303_n388#
+ a_n465_n388# a_447_n300# a_399_322# a_159_n300# a_111_n388# a_15_322# a_n273_n388#
+ a_255_n300# a_n611_n474# a_351_n300# a_207_322# a_n417_n300# a_n129_n300# a_n81_n388#
+ a_63_n300# a_n177_322# a_n225_n300# a_n321_n300#
X0 a_255_n300# a_207_322# a_159_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X1 a_n321_n300# a_n369_322# a_n417_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X2 a_159_n300# a_111_n388# a_63_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X3 a_n225_n300# a_n273_n388# a_n321_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X4 a_447_n300# a_399_322# a_351_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X5 a_63_n300# a_15_322# a_n33_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X6 a_n129_n300# a_n177_322# a_n225_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X7 a_n417_n300# a_n465_n388# a_n509_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X8 a_n33_n300# a_n81_n388# a_n129_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X9 a_351_n300# a_303_n388# a_255_n300# a_n611_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_VC5YSW a_63_n800# a_n81_831# a_n225_n800# a_15_n897#
+ a_n177_n897# a_n561_n897# a_927_n800# a_879_831# a_n273_831# a_n321_n800# a_639_n800#
+ a_735_n800# a_n33_n800# a_n465_831# a_n897_n800# a_831_n800# a_447_n800# a_783_n897#
+ a_399_n897# a_543_n800# a_159_n800# a_n609_n800# a_n945_n897# a_n657_831# a_495_831#
+ a_255_n800# a_n705_n800# a_111_831# a_591_n897# a_207_n897# w_n1127_n1019# a_351_n800#
+ a_n417_n800# a_n801_n800# a_n753_n897# a_n849_831# a_n369_n897# a_687_831# a_303_831#
+ a_n129_n800# a_n513_n800# a_n989_n800#
X0 a_n33_n800# a_n81_831# a_n129_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1 a_351_n800# a_303_831# a_255_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2 a_n609_n800# a_n657_831# a_n705_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3 a_927_n800# a_879_831# a_831_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X4 a_n897_n800# a_n945_n897# a_n989_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
X5 a_255_n800# a_207_n897# a_159_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6 a_n321_n800# a_n369_n897# a_n417_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X7 a_543_n800# a_495_831# a_447_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8 a_831_n800# a_783_n897# a_735_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X9 a_159_n800# a_111_831# a_63_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X10 a_n225_n800# a_n273_831# a_n321_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X11 a_447_n800# a_399_n897# a_351_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X12 a_n513_n800# a_n561_n897# a_n609_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X13 a_63_n800# a_15_n897# a_n33_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X14 a_735_n800# a_687_831# a_639_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X15 a_n801_n800# a_n849_831# a_n897_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X16 a_n129_n800# a_n177_n897# a_n225_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X17 a_n417_n800# a_n465_831# a_n513_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X18 a_639_n800# a_591_n897# a_543_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X19 a_n705_n800# a_n753_n897# a_n801_n800# w_n1127_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_Z85QYA a_n753_n388# a_n849_322# a_735_n300# a_n33_n300#
+ a_n369_n388# a_687_322# a_303_322# a_n897_n300# a_831_n300# a_447_n300# a_15_n388#
+ a_n81_322# a_n177_n388# a_n561_n388# a_543_n300# a_159_n300# a_n609_n300# a_879_322#
+ a_n273_322# a_255_n300# a_n705_n300# a_351_n300# a_n801_n300# a_n417_n300# a_n465_322#
+ a_n513_n300# a_n989_n300# a_n129_n300# a_783_n388# a_399_n388# a_63_n300# a_n225_n300#
+ a_n657_322# a_n945_n388# a_927_n300# a_n1091_n474# a_495_322# a_n321_n300# a_591_n388#
+ a_111_322# a_639_n300# a_207_n388#
X0 a_n897_n300# a_n945_n388# a_n989_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X1 a_927_n300# a_879_322# a_831_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X2 a_255_n300# a_207_n388# a_159_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X3 a_n321_n300# a_n369_n388# a_n417_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X4 a_543_n300# a_495_322# a_447_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X5 a_831_n300# a_783_n388# a_735_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X6 a_159_n300# a_111_322# a_63_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X7 a_n225_n300# a_n273_322# a_n321_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X8 a_447_n300# a_399_n388# a_351_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X9 a_n513_n300# a_n561_n388# a_n609_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X10 a_63_n300# a_15_n388# a_n33_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X11 a_735_n300# a_687_322# a_639_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X12 a_n801_n300# a_n849_322# a_n897_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X13 a_n129_n300# a_n177_n388# a_n225_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X14 a_n417_n300# a_n465_322# a_n513_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X15 a_639_n300# a_591_n388# a_543_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X16 a_n705_n300# a_n753_n388# a_n801_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X17 a_n33_n300# a_n81_322# a_n129_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X18 a_351_n300# a_303_322# a_255_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X19 a_n609_n300# a_n657_322# a_n705_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
.ends

.subckt sky130_fd_pr__nfet_01v8_PPAFLS a_n753_n388# a_n849_322# a_735_n300# a_n33_n300#
+ a_n369_n388# a_687_322# a_303_322# a_n897_n300# a_831_n300# a_447_n300# a_15_n388#
+ a_n81_322# a_n177_n388# a_n561_n388# a_543_n300# a_159_n300# a_n609_n300# a_879_322#
+ a_n273_322# a_255_n300# a_n705_n300# a_351_n300# a_n801_n300# a_n417_n300# a_n465_322#
+ a_n513_n300# a_n989_n300# a_n129_n300# a_783_n388# a_399_n388# a_63_n300# a_n225_n300#
+ a_n657_322# a_n945_n388# a_927_n300# a_n1091_n474# a_495_322# a_n321_n300# a_591_n388#
+ a_111_322# a_639_n300# a_207_n388#
X0 a_n897_n300# a_n945_n388# a_n989_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X1 a_927_n300# a_879_322# a_831_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X2 a_255_n300# a_207_n388# a_159_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X3 a_n321_n300# a_n369_n388# a_n417_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X4 a_543_n300# a_495_322# a_447_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X5 a_831_n300# a_783_n388# a_735_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X6 a_159_n300# a_111_322# a_63_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X7 a_n225_n300# a_n273_322# a_n321_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X8 a_447_n300# a_399_n388# a_351_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X9 a_n513_n300# a_n561_n388# a_n609_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X10 a_63_n300# a_15_n388# a_n33_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X11 a_735_n300# a_687_322# a_639_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X12 a_n801_n300# a_n849_322# a_n897_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X13 a_n129_n300# a_n177_n388# a_n225_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X14 a_n417_n300# a_n465_322# a_n513_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X15 a_639_n300# a_591_n388# a_543_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X16 a_n705_n300# a_n753_n388# a_n801_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X17 a_n33_n300# a_n81_322# a_n129_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X18 a_351_n300# a_303_322# a_255_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X19 a_n609_n300# a_n657_322# a_n705_n300# a_n1091_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
.ends

.subckt vco vdd out vctrl vss
XXM12 w_8958_n708# w_8958_n708# w_8958_n708# out m1_6574_n1254# m1_6574_n1254# out
+ out m1_6574_n1254# out m1_6574_n1254# m1_6574_n1254# m1_6574_n1254# w_8958_n708#
+ m1_6574_n1254# m1_6574_n1254# m1_6574_n1254# w_8958_n708# w_8958_n708# w_8958_n708#
+ m1_6574_n1254# m1_6574_n1254# m1_6574_n1254# out out m1_6574_n1254# m1_6574_n1254#
+ w_8958_n708# w_8958_n708# m1_6574_n1254# w_8958_n708# w_8958_n708# m1_6574_n1254#
+ m1_6574_n1254# m1_6574_n1254# out m1_6574_n1254# out m1_6574_n1254# out out m1_6574_n1254#
+ m1_6574_n1254# w_8958_n708# w_8958_n708# m1_6574_n1254# m1_6574_n1254# w_8958_n708#
+ w_8958_n708# m1_6574_n1254# out out out m1_6574_n1254# out out m1_6574_n1254# m1_6574_n1254#
+ w_8958_n708# w_8958_n708# m1_6574_n1254# m1_6574_n1254# sky130_fd_pr__pfet_01v8_VC56GX
XXM14 m1_6574_n1254# m1_9090_n2156# m1_9090_n2156# m1_6574_n1254# m1_6574_n1254# out
+ m1_6574_n1254# out m1_6574_n1254# m1_6574_n1254# out out m1_9090_n2156# m1_6574_n1254#
+ m1_6574_n1254# m1_9090_n2156# m1_9090_n2156# m1_9090_n2156# m1_6574_n1254# m1_6574_n1254#
+ m1_6574_n1254# m1_6574_n1254# m1_6574_n1254# m1_6574_n1254# m1_6574_n1254# out out
+ out m1_6574_n1254# m1_6574_n1254# vss m1_9090_n2156# m1_9090_n2156# m1_6574_n1254#
+ m1_9090_n2156# m1_6574_n1254# m1_6574_n1254# m1_9090_n2156# m1_9090_n2156# m1_6574_n1254#
+ out out m1_6574_n1254# m1_6574_n1254# m1_6574_n1254# out out out m1_6574_n1254#
+ m1_6574_n1254# m1_9090_n2156# m1_6574_n1254# m1_9090_n2156# m1_9090_n2156# m1_9090_n2156#
+ m1_6574_n1254# out m1_6574_n1254# m1_6574_n1254# out out out sky130_fd_pr__nfet_01v8_UBPJLS
XXM13 vctrl vss vss vctrl vctrl m1_9090_n2156# vctrl m1_9090_n2156# vctrl vctrl m1_9090_n2156#
+ m1_9090_n2156# vss vctrl vctrl vss vss vss vctrl vctrl vctrl vctrl vctrl vctrl vctrl
+ m1_9090_n2156# m1_9090_n2156# m1_9090_n2156# vctrl vctrl vss vss vss vctrl vss vctrl
+ vctrl vss vss vctrl m1_9090_n2156# m1_9090_n2156# vctrl vctrl vctrl m1_9090_n2156#
+ m1_9090_n2156# m1_9090_n2156# vctrl vctrl vss vctrl vss vss vss vctrl m1_9090_n2156#
+ vctrl vctrl m1_9090_n2156# m1_9090_n2156# m1_9090_n2156# sky130_fd_pr__nfet_01v8_CDSMYA
XXM1 vss vss vctrl vctrl m1_3928_n926# vss vctrl m1_3928_n926# m1_3928_n926# vss vctrl
+ vctrl sky130_fd_pr__nfet_01v8_42S873
XXM2 vdd m1_3928_n926# m1_3928_n926# vdd m1_3928_n926# vdd m1_3928_n926# m1_3928_n926#
+ vdd m1_3928_n926# m1_3928_n926# m1_3928_n926# sky130_fd_pr__pfet_01v8_UYM7GH
XXM3 vdd w_4930_1018# vdd m1_3928_n926# m1_3928_n926# w_4930_1018# m1_3928_n926# m1_3928_n926#
+ m1_3928_n926# vdd w_4930_1018# w_4930_1018# m1_3928_n926# m1_3928_n926# vdd w_4930_1018#
+ m1_3928_n926# vdd vdd m1_3928_n926# w_4930_1018# m1_3928_n926# sky130_fd_pr__pfet_01v8_VC5S4W
XXM4 w_4930_1018# w_4930_1018# m1_5022_n1250# out out w_4930_1018# out out out m1_5022_n1250#
+ w_4930_1018# w_4930_1018# out out m1_5022_n1250# w_4930_1018# out m1_5022_n1250#
+ m1_5022_n1250# out w_4930_1018# out sky130_fd_pr__pfet_01v8_VC5S4W
XXM5 vctrl vss m1_5024_n2164# vctrl vctrl m1_5024_n2164# vctrl vss vctrl vctrl vctrl
+ m1_5024_n2164# vss vss vctrl vss m1_5024_n2164# vctrl m1_5024_n2164# vctrl vss m1_5024_n2164#
+ sky130_fd_pr__nfet_01v8_JT8PYA
XXM6 out m1_5024_n2164# m1_5022_n1250# out out m1_5022_n1250# out m1_5024_n2164# out
+ out out m1_5022_n1250# vss m1_5024_n2164# out m1_5024_n2164# m1_5022_n1250# out
+ m1_5022_n1250# out m1_5024_n2164# m1_5022_n1250# sky130_fd_pr__nfet_01v8_JLF2PR
XXM7 vdd m1_3928_n926# m1_6572_874# m1_3928_n926# m1_3928_n926# m1_3928_n926# m1_6572_874#
+ m1_3928_n926# m1_3928_n926# vdd vdd m1_6572_874# m1_6572_874# m1_3928_n926# vdd
+ vdd vdd m1_3928_n926# m1_3928_n926# m1_6572_874# m1_6572_874# m1_6572_874# m1_3928_n926#
+ m1_3928_n926# m1_3928_n926# vdd vdd m1_3928_n926# m1_3928_n926# m1_3928_n926# vdd
+ m1_6572_874# m1_6572_874# m1_6572_874# m1_3928_n926# m1_3928_n926# m1_3928_n926#
+ m1_3928_n926# m1_3928_n926# vdd vdd m1_6572_874# sky130_fd_pr__pfet_01v8_VC5YSW
XXM8 m1_6574_n1254# m1_5022_n1250# m1_6572_874# m1_5022_n1250# m1_5022_n1250# m1_5022_n1250#
+ m1_6572_874# m1_5022_n1250# m1_5022_n1250# m1_6574_n1254# m1_6574_n1254# m1_6572_874#
+ m1_6572_874# m1_5022_n1250# m1_6574_n1254# m1_6574_n1254# m1_6574_n1254# m1_5022_n1250#
+ m1_5022_n1250# m1_6572_874# m1_6572_874# m1_6572_874# m1_5022_n1250# m1_5022_n1250#
+ m1_5022_n1250# m1_6574_n1254# m1_6574_n1254# m1_5022_n1250# m1_5022_n1250# m1_5022_n1250#
+ m1_6572_874# m1_6572_874# m1_6572_874# m1_6572_874# m1_5022_n1250# m1_5022_n1250#
+ m1_5022_n1250# m1_5022_n1250# m1_5022_n1250# m1_6574_n1254# m1_6574_n1254# m1_6572_874#
+ sky130_fd_pr__pfet_01v8_VC5YSW
XXM9 vctrl vctrl m1_6574_n2166# m1_6574_n2166# vctrl vctrl vctrl vss vss vss vctrl
+ vctrl vctrl vctrl m1_6574_n2166# m1_6574_n2166# m1_6574_n2166# vctrl vctrl vss vss
+ m1_6574_n2166# m1_6574_n2166# m1_6574_n2166# vctrl vss m1_6574_n2166# vss vctrl
+ vctrl vss m1_6574_n2166# vctrl vctrl m1_6574_n2166# vss vctrl vss vctrl vctrl vss
+ vctrl sky130_fd_pr__nfet_01v8_Z85QYA
XXM10 m1_5022_n1250# m1_5022_n1250# m1_6574_n1254# m1_6574_n1254# m1_5022_n1250# m1_5022_n1250#
+ m1_5022_n1250# m1_6574_n2166# m1_6574_n2166# m1_6574_n2166# m1_5022_n1250# m1_5022_n1250#
+ m1_5022_n1250# m1_5022_n1250# m1_6574_n1254# m1_6574_n1254# m1_6574_n1254# m1_5022_n1250#
+ m1_5022_n1250# m1_6574_n2166# m1_6574_n2166# m1_6574_n1254# m1_6574_n1254# m1_6574_n1254#
+ m1_5022_n1250# m1_6574_n2166# m1_6574_n1254# m1_6574_n2166# m1_5022_n1250# m1_5022_n1250#
+ m1_6574_n2166# m1_6574_n1254# m1_5022_n1250# m1_5022_n1250# m1_6574_n1254# vss m1_5022_n1250#
+ m1_6574_n2166# m1_5022_n1250# m1_5022_n1250# m1_6574_n2166# m1_5022_n1250# sky130_fd_pr__nfet_01v8_PPAFLS
XXM11 w_8958_n708# w_8958_n708# w_8958_n708# vdd m1_3928_n926# m1_3928_n926# vdd vdd
+ m1_3928_n926# vdd m1_3928_n926# m1_3928_n926# m1_3928_n926# w_8958_n708# m1_3928_n926#
+ m1_3928_n926# m1_3928_n926# w_8958_n708# w_8958_n708# w_8958_n708# m1_3928_n926#
+ m1_3928_n926# m1_3928_n926# vdd vdd m1_3928_n926# m1_3928_n926# w_8958_n708# w_8958_n708#
+ m1_3928_n926# w_8958_n708# w_8958_n708# m1_3928_n926# m1_3928_n926# m1_3928_n926#
+ vdd m1_3928_n926# vdd m1_3928_n926# vdd vdd m1_3928_n926# m1_3928_n926# w_8958_n708#
+ w_8958_n708# m1_3928_n926# m1_3928_n926# w_8958_n708# vdd m1_3928_n926# vdd vdd
+ vdd m1_3928_n926# vdd vdd m1_3928_n926# m1_3928_n926# w_8958_n708# w_8958_n708#
+ m1_3928_n926# m1_3928_n926# sky130_fd_pr__pfet_01v8_VC56GX
.ends

