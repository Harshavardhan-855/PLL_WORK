magic
tech sky130A
magscale 1 2
timestamp 1709895641
<< nwell >>
rect 3997 101 4202 399
rect 3982 -458 4309 -304
rect 3982 -602 4310 -458
rect 4000 -626 4310 -602
rect 3988 -1304 4279 -1006
rect 3988 -1306 4078 -1304
<< pwell >>
rect 3958 -160 4094 22
rect 3962 -866 4102 -682
rect 3950 -1568 4112 -1384
<< psubdiff >>
rect 3988 -12 4062 12
rect 3988 -152 4062 -128
rect 3992 -708 4062 -684
rect 3992 -854 4062 -830
rect 3994 -1404 4060 -1380
rect 3994 -1568 4060 -1544
<< nsubdiff >>
rect 3997 329 4022 363
rect 4106 329 4166 363
rect 4132 303 4166 329
rect 4132 171 4166 197
rect 3997 137 4022 171
rect 4106 137 4166 171
rect 4104 -378 4129 -344
rect 4213 -378 4273 -344
rect 4239 -404 4273 -378
rect 4239 -536 4273 -510
rect 4104 -570 4129 -536
rect 4213 -570 4273 -536
rect 4074 -1076 4099 -1042
rect 4183 -1076 4243 -1042
rect 4209 -1102 4243 -1076
rect 4209 -1234 4243 -1208
rect 4074 -1268 4099 -1234
rect 4183 -1268 4243 -1234
<< psubdiffcont >>
rect 3988 -128 4062 -12
rect 3992 -830 4062 -708
rect 3994 -1544 4060 -1404
<< nsubdiffcont >>
rect 4022 329 4106 363
rect 4132 197 4166 303
rect 4022 137 4106 171
rect 4129 -378 4213 -344
rect 4239 -510 4273 -404
rect 4129 -570 4213 -536
rect 4099 -1076 4183 -1042
rect 4209 -1208 4243 -1102
rect 4099 -1268 4183 -1234
<< locali >>
rect 3940 326 4022 380
rect 4106 329 4166 363
rect 4132 303 4166 329
rect 4132 171 4166 197
rect 3997 137 4022 171
rect 4106 137 4166 171
rect 1744 36 2094 72
rect 3988 -12 4062 4
rect 3988 -164 4062 -128
rect 1936 -198 2172 -164
rect 3940 -180 4062 -164
rect 3958 -198 4062 -180
rect 1938 -870 1980 -198
rect 3944 -344 4036 -324
rect 3944 -358 4129 -344
rect 4002 -378 4129 -358
rect 4213 -378 4273 -344
rect 4239 -404 4273 -378
rect 4239 -536 4273 -510
rect 4104 -570 4129 -536
rect 4213 -570 4273 -536
rect 3992 -708 4062 -692
rect 3992 -846 4062 -830
rect 1938 -880 2174 -870
rect 1936 -904 2174 -880
rect 3942 -904 4060 -846
rect 1936 -1570 1986 -904
rect 3918 -1028 4074 -1024
rect 3950 -1042 4074 -1028
rect 3950 -1058 4099 -1042
rect 3996 -1076 4099 -1058
rect 4183 -1076 4243 -1042
rect 4209 -1102 4243 -1076
rect 4209 -1234 4243 -1208
rect 4074 -1268 4099 -1234
rect 4183 -1268 4243 -1234
rect 3994 -1404 4060 -1388
rect 3410 -1512 3456 -1504
rect 3994 -1566 4060 -1544
rect 1762 -1606 2164 -1570
rect 3928 -1604 4060 -1566
rect 1936 -1608 1986 -1606
<< viali >>
rect 3798 120 3836 158
rect 1708 36 1744 72
rect 2304 22 2348 62
rect 3414 -96 3460 -50
rect 3800 -580 3844 -540
rect 2052 -688 2108 -632
rect 2308 -696 2360 -650
rect 3424 -802 3470 -756
rect 1720 -1608 1762 -1568
rect 3790 -1284 3836 -1242
rect 2038 -1388 2102 -1334
rect 2302 -1384 2344 -1344
rect 3410 -1504 3456 -1466
<< metal1 >>
rect 1588 314 2056 410
rect 1588 210 1788 314
rect 1592 72 1792 82
rect 1592 36 1708 72
rect 1744 36 1792 72
rect 1592 -118 1792 36
rect 1868 -298 1908 314
rect 3786 158 3848 164
rect 3786 120 3798 158
rect 3836 120 3848 158
rect 3786 114 3848 120
rect 2290 70 2348 74
rect 3786 70 3846 114
rect 2290 68 3846 70
rect 2290 16 2300 68
rect 2358 16 3846 68
rect 2294 14 3846 16
rect 2348 12 2376 14
rect 4138 -34 4338 38
rect 3396 -102 3406 -42
rect 3468 -102 3478 -42
rect 4138 -98 4174 -34
rect 4228 -98 4338 -34
rect 4138 -162 4338 -98
rect 1868 -304 1912 -298
rect 1868 -384 2126 -304
rect 1868 -1006 1912 -384
rect 3788 -540 3856 -534
rect 3788 -580 3800 -540
rect 3844 -580 3856 -540
rect 3788 -586 3856 -580
rect 2028 -694 2038 -622
rect 2102 -626 2112 -622
rect 2102 -632 2120 -626
rect 2108 -688 2120 -632
rect 2306 -634 2360 -630
rect 3802 -634 3854 -586
rect 2306 -642 3856 -634
rect 2102 -694 2120 -688
rect 2292 -694 2302 -642
rect 2366 -676 3856 -642
rect 2366 -694 3708 -676
rect 2296 -696 2308 -694
rect 2360 -696 3708 -694
rect 2296 -702 3708 -696
rect 4148 -740 4348 -678
rect 3408 -808 3418 -750
rect 3476 -808 3486 -750
rect 4148 -816 4188 -740
rect 4244 -816 4348 -740
rect 4148 -878 4348 -816
rect 1870 -1008 1912 -1006
rect 1870 -1088 2146 -1008
rect 3778 -1242 3848 -1236
rect 3778 -1284 3790 -1242
rect 3836 -1284 3848 -1242
rect 3778 -1290 3848 -1284
rect 2020 -1394 2030 -1326
rect 2098 -1328 2108 -1326
rect 2098 -1334 2114 -1328
rect 2102 -1388 2114 -1334
rect 2290 -1340 2356 -1338
rect 2098 -1394 2114 -1388
rect 2288 -1342 3668 -1340
rect 3790 -1342 3836 -1290
rect 2288 -1344 3838 -1342
rect 2288 -1384 2302 -1344
rect 2344 -1384 3838 -1344
rect 2288 -1390 3838 -1384
rect 2288 -1392 3668 -1390
rect 1590 -1568 1792 -1432
rect 4158 -1446 4358 -1382
rect 3398 -1458 3468 -1452
rect 3388 -1510 3398 -1458
rect 3462 -1510 3472 -1458
rect 4158 -1510 4196 -1446
rect 4260 -1510 4358 -1446
rect 1590 -1608 1720 -1568
rect 1762 -1608 1792 -1568
rect 4158 -1582 4358 -1510
rect 1590 -1634 1792 -1608
<< via1 >>
rect 2300 62 2358 68
rect 2300 22 2304 62
rect 2304 22 2348 62
rect 2348 22 2358 62
rect 2300 16 2358 22
rect 3406 -50 3468 -42
rect 3406 -96 3414 -50
rect 3414 -96 3460 -50
rect 3460 -96 3468 -50
rect 3406 -102 3468 -96
rect 4174 -98 4228 -34
rect 2038 -632 2102 -622
rect 2038 -688 2052 -632
rect 2052 -688 2102 -632
rect 2038 -694 2102 -688
rect 2302 -650 2366 -642
rect 2302 -694 2308 -650
rect 2308 -694 2360 -650
rect 2360 -694 2366 -650
rect 3418 -756 3476 -750
rect 3418 -802 3424 -756
rect 3424 -802 3470 -756
rect 3470 -802 3476 -756
rect 3418 -808 3476 -802
rect 4188 -816 4244 -740
rect 2030 -1334 2098 -1326
rect 2030 -1388 2038 -1334
rect 2038 -1388 2098 -1334
rect 2030 -1394 2098 -1388
rect 3398 -1466 3462 -1458
rect 3398 -1504 3410 -1466
rect 3410 -1504 3456 -1466
rect 3456 -1504 3462 -1466
rect 3398 -1510 3462 -1504
rect 4196 -1510 4260 -1446
<< metal2 >>
rect 2300 68 2358 78
rect 2358 16 2360 48
rect 2300 -244 2360 16
rect 3406 -42 3468 -32
rect 4174 -34 4228 -24
rect 3468 -92 4174 -44
rect 3406 -112 3468 -102
rect 4174 -108 4228 -98
rect 2040 -294 2360 -244
rect 2040 -612 2102 -294
rect 2038 -622 2102 -612
rect 2038 -704 2102 -694
rect 2302 -642 2366 -632
rect 2302 -704 2366 -694
rect 2306 -948 2364 -704
rect 4188 -740 4244 -730
rect 3418 -750 3476 -740
rect 4090 -752 4188 -750
rect 3476 -808 4188 -752
rect 3418 -818 3476 -808
rect 4188 -826 4244 -816
rect 2044 -988 2364 -948
rect 2044 -1316 2088 -988
rect 2030 -1326 2098 -1316
rect 2030 -1404 2098 -1394
rect 4196 -1446 4260 -1436
rect 3398 -1458 4196 -1446
rect 3462 -1510 4196 -1458
rect 4260 -1510 4262 -1446
rect 3398 -1520 3462 -1510
rect 4196 -1520 4260 -1510
use sky130_fd_sc_hd__dfxbp_2  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1705271942
transform 1 0 2032 0 1 -886
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_2  x2
timestamp 1705271942
transform 1 0 2020 0 1 -1588
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_2  x3
timestamp 1705271942
transform 1 0 2028 0 1 -182
box -38 -48 1970 592
<< labels >>
flabel metal1 4138 -162 4338 38 0 FreeSans 256 0 0 0 out_a
port 1 nsew
flabel metal1 4148 -878 4348 -678 0 FreeSans 256 0 0 0 out_b
port 2 nsew
flabel metal1 4158 -1582 4358 -1382 0 FreeSans 256 0 0 0 out_c
port 3 nsew
flabel metal1 1590 -1634 1790 -1434 0 FreeSans 256 0 0 0 vss
port 5 nsew
flabel metal1 1588 210 1788 410 0 FreeSans 256 0 0 0 vdd
port 4 nsew
flabel metal1 1592 -118 1792 82 0 FreeSans 256 0 0 0 clock
port 0 nsew
<< end >>
