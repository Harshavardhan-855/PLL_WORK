magic
tech sky130A
magscale 1 2
timestamp 1709641130
<< nwell >>
rect 2546 416 3364 422
rect 2524 300 3364 416
rect 3306 168 3364 300
<< locali >>
rect 2440 1494 2594 1528
rect 3072 1382 3110 1526
rect 3906 1380 3954 1528
rect 4202 1236 4324 1296
rect 4392 542 4426 666
rect 4398 192 4432 326
rect 3822 -24 3858 120
rect 3818 -374 3854 -244
rect 4190 -696 4298 -658
rect 4282 -920 4700 -872
<< viali >>
rect 2404 1494 2440 1528
rect 4700 -920 4750 -868
<< metal1 >>
rect 2324 1528 2524 1562
rect 2324 1494 2404 1528
rect 2440 1494 2524 1528
rect 2324 1362 2524 1494
rect 3184 1486 4422 1542
rect 2736 1378 2746 1430
rect 2850 1378 2860 1430
rect 3184 1376 3242 1486
rect 4358 1446 4422 1486
rect 2642 596 2704 1374
rect 3030 1254 3040 1306
rect 3144 1254 3154 1306
rect 2736 1138 2746 1190
rect 2850 1138 2860 1190
rect 3026 1018 3036 1070
rect 3140 1018 3150 1070
rect 2732 900 2742 952
rect 2846 900 2856 952
rect 3028 780 3038 832
rect 3142 780 3152 832
rect 2736 662 2746 714
rect 2850 662 2860 714
rect 3182 596 3244 1376
rect 3568 1374 3578 1426
rect 3682 1374 3692 1426
rect 4358 1390 4662 1446
rect 3024 540 3034 592
rect 3138 540 3148 592
rect 3108 508 3142 540
rect 2320 432 2520 506
rect 3108 498 3228 508
rect 3108 470 3230 498
rect 3122 468 3230 470
rect 2320 354 2380 432
rect 2454 354 2520 432
rect 2320 306 2520 354
rect 3194 110 3230 468
rect 3462 418 3526 1370
rect 3822 1254 3832 1306
rect 3954 1254 3964 1306
rect 3568 1136 3578 1188
rect 3682 1136 3692 1188
rect 3822 1018 3832 1070
rect 3954 1018 3964 1070
rect 3568 900 3578 952
rect 3682 900 3692 952
rect 3822 782 3832 834
rect 3954 782 3964 834
rect 3568 664 3578 716
rect 3682 664 3692 716
rect 3810 546 3820 598
rect 3954 546 3964 598
rect 3568 428 3578 480
rect 3682 428 3692 480
rect 3448 358 3458 418
rect 3516 358 3526 418
rect 3462 354 3526 358
rect 3812 306 3822 364
rect 3958 306 3968 364
rect 4004 362 4068 1378
rect 4294 1200 4304 1336
rect 4360 1200 4370 1336
rect 4532 1200 4542 1336
rect 4598 1200 4608 1336
rect 4412 958 4422 1096
rect 4478 958 4488 1096
rect 4650 958 4660 1096
rect 4716 958 4726 1096
rect 4656 902 4726 958
rect 4598 900 4726 902
rect 4358 844 4726 900
rect 4466 762 4532 844
rect 4456 678 4466 762
rect 4530 678 4540 762
rect 4304 408 4364 534
rect 4394 414 4404 474
rect 4592 414 4600 474
rect 4632 411 4692 534
rect 4152 350 4364 408
rect 4152 348 4336 350
rect 3166 96 3230 110
rect 3130 34 3230 96
rect 2324 -130 2524 -60
rect 2324 -190 2398 -130
rect 2452 -190 2524 -130
rect 2324 -260 2524 -190
rect 2610 -86 2702 -34
rect 2610 -94 2674 -86
rect 2610 -346 2658 -94
rect 2710 -190 2720 -132
rect 2782 -190 2792 -132
rect 3730 -218 3788 -30
rect 4152 -44 4192 348
rect 4052 -84 4192 -44
rect 3822 -152 3832 -98
rect 4006 -104 4016 -98
rect 4052 -104 4110 -84
rect 4006 -142 4110 -104
rect 4006 -152 4016 -142
rect 4052 -166 4110 -142
rect 4052 -206 4160 -166
rect 2592 -412 2602 -346
rect 2664 -412 2674 -346
rect 2320 -516 2520 -442
rect 2320 -574 2386 -516
rect 2444 -574 2520 -516
rect 2320 -642 2520 -574
rect 2610 -600 2658 -412
rect 2706 -574 2716 -514
rect 2774 -574 2784 -514
rect 4098 -520 4160 -206
rect 4650 -342 4850 -270
rect 4650 -416 4688 -342
rect 4760 -416 4850 -342
rect 4650 -470 4850 -416
rect 4094 -572 4162 -520
rect 2610 -616 2680 -600
rect 2610 -668 2706 -616
rect 3726 -732 4082 -678
rect 4086 -836 4158 -778
rect 4658 -868 4858 -816
rect 4658 -920 4700 -868
rect 4750 -920 4858 -868
rect 4658 -1016 4858 -920
<< via1 >>
rect 2746 1378 2850 1430
rect 3040 1254 3144 1306
rect 2746 1138 2850 1190
rect 3036 1018 3140 1070
rect 2742 900 2846 952
rect 3038 780 3142 832
rect 2746 662 2850 714
rect 3578 1374 3682 1426
rect 3034 540 3138 592
rect 2380 354 2454 432
rect 3832 1254 3954 1306
rect 3578 1136 3682 1188
rect 3832 1018 3954 1070
rect 3578 900 3682 952
rect 3832 782 3954 834
rect 3578 664 3682 716
rect 3820 546 3954 598
rect 3578 428 3682 480
rect 3458 358 3516 418
rect 3822 306 3958 364
rect 4304 1200 4360 1336
rect 4542 1200 4598 1336
rect 4422 958 4478 1096
rect 4660 958 4716 1096
rect 4466 678 4530 762
rect 4404 414 4592 474
rect 2398 -190 2452 -130
rect 2720 -190 2782 -132
rect 3832 -152 4006 -98
rect 2602 -412 2664 -346
rect 2386 -574 2444 -516
rect 2716 -574 2774 -514
rect 4688 -416 4760 -342
<< metal2 >>
rect 2746 1430 2850 1440
rect 3578 1432 3682 1436
rect 2738 1378 2746 1430
rect 2850 1378 2852 1430
rect 2738 1190 2852 1378
rect 3572 1426 3682 1432
rect 3572 1374 3578 1426
rect 3572 1364 3682 1374
rect 3040 1308 3144 1316
rect 3040 1306 3146 1308
rect 3144 1254 3146 1306
rect 3040 1244 3146 1254
rect 2738 1138 2746 1190
rect 2850 1138 2852 1190
rect 2738 952 2852 1138
rect 3044 1080 3146 1244
rect 3036 1070 3146 1080
rect 3140 1018 3146 1070
rect 3036 1008 3146 1018
rect 2738 900 2742 952
rect 2846 900 2852 952
rect 2738 714 2852 900
rect 3044 842 3146 1008
rect 3038 832 3146 842
rect 3142 780 3146 832
rect 3038 770 3146 780
rect 2738 662 2746 714
rect 2850 662 2852 714
rect 2746 652 2850 662
rect 3044 602 3146 770
rect 3034 592 3146 602
rect 3138 540 3146 592
rect 3034 538 3146 540
rect 3572 1198 3680 1364
rect 4304 1338 4360 1346
rect 4542 1338 4598 1346
rect 4302 1336 4600 1338
rect 3832 1308 3954 1316
rect 3832 1306 3958 1308
rect 3954 1254 3958 1306
rect 3572 1188 3682 1198
rect 3572 1136 3578 1188
rect 3572 1126 3682 1136
rect 3572 962 3680 1126
rect 3832 1070 3958 1254
rect 4302 1200 4304 1336
rect 4360 1200 4542 1336
rect 4598 1200 4600 1336
rect 4304 1190 4360 1200
rect 4542 1190 4598 1200
rect 4422 1098 4478 1106
rect 4660 1098 4716 1106
rect 3954 1018 3958 1070
rect 3572 952 3682 962
rect 3572 900 3578 952
rect 3572 890 3682 900
rect 3572 726 3680 890
rect 3832 834 3958 1018
rect 4416 1096 4718 1098
rect 4416 958 4422 1096
rect 4478 958 4660 1096
rect 4716 958 4718 1096
rect 4416 956 4718 958
rect 4422 948 4478 956
rect 4660 948 4716 956
rect 3954 782 3958 834
rect 3572 716 3682 726
rect 3572 664 3578 716
rect 3572 654 3682 664
rect 3034 530 3138 538
rect 3572 490 3680 654
rect 3832 608 3958 782
rect 3820 598 3958 608
rect 3954 546 3958 598
rect 3820 536 3958 546
rect 3572 480 3682 490
rect 2380 432 2454 442
rect 3572 428 3578 480
rect 3458 420 3516 428
rect 2454 418 3516 420
rect 2454 358 3458 418
rect 3572 418 3682 428
rect 3572 416 3680 418
rect 3832 374 3958 536
rect 4466 762 4530 772
rect 4466 668 4530 678
rect 4466 484 4528 668
rect 4404 474 4592 484
rect 4404 404 4592 414
rect 2454 354 3516 358
rect 2380 344 2454 354
rect 3458 348 3516 354
rect 3822 364 3958 374
rect 3822 296 3958 306
rect 3866 -88 3942 296
rect 3832 -98 4006 -88
rect 2398 -130 2452 -120
rect 2720 -132 2782 -122
rect 2452 -188 2720 -134
rect 2398 -200 2452 -190
rect 3832 -162 4006 -152
rect 2720 -200 2782 -190
rect 2602 -342 2664 -336
rect 4688 -342 4760 -332
rect 2598 -346 4688 -342
rect 2598 -412 2602 -346
rect 2664 -412 4688 -346
rect 2598 -416 4688 -412
rect 2602 -422 2664 -416
rect 4688 -426 4760 -416
rect 2386 -516 2444 -506
rect 2716 -514 2774 -504
rect 2444 -572 2716 -516
rect 2386 -584 2444 -574
rect 2716 -584 2774 -574
use sky130_fd_pr__pfet_01v8_6QKSWZ  XM1
timestamp 1709561889
transform 1 0 4510 0 1 1147
box -344 -419 344 419
use sky130_fd_pr__nfet_01v8_8LLW3F  XM2
timestamp 1709561889
transform 0 1 4496 -1 0 441
box -285 -310 285 310
use sky130_fd_pr__nfet_01v8_8LLW3F  XM3
timestamp 1709561889
transform 0 -1 3920 1 0 -125
box -285 -310 285 310
use sky130_fd_pr__pfet_01v8_6Q3TWZ  XM4
timestamp 1709561889
transform 0 1 2943 -1 0 984
box -580 -419 580 419
use sky130_fd_pr__nfet_01v8_8YFQNF  XM5
timestamp 1709561889
transform -1 0 4126 0 -1 -676
box -226 -280 226 280
use sky130_fd_pr__pfet_01v8_GJYSVV  XM6
timestamp 1709561889
transform 1 0 2920 0 1 7
box -396 -319 396 319
use sky130_fd_pr__nfet_01v8_U4BYG2  XM7
timestamp 1709561889
transform 1 0 3216 0 1 -704
box -696 -310 696 310
use sky130_fd_pr__pfet_01v8_6QBZWZ  XM8
timestamp 1709561889
transform 0 1 3765 1 0 866
box -698 -419 698 419
<< labels >>
flabel metal1 2320 306 2520 506 0 FreeSans 256 0 0 0 cp_bias
port 1 nsew
flabel metal1 2324 -260 2524 -60 0 FreeSans 256 0 0 0 qa
port 2 nsew
flabel metal1 2320 -642 2520 -442 0 FreeSans 256 0 0 0 qb
port 4 nsew
flabel metal1 4650 -470 4850 -270 0 FreeSans 256 0 0 0 cp_out
port 3 nsew
flabel metal1 4658 -1016 4858 -816 0 FreeSans 256 0 0 0 vss
port 5 nsew
flabel metal1 2324 1362 2524 1562 0 FreeSans 256 0 0 0 vdd
port 0 nsew
<< end >>
