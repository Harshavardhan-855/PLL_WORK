magic
tech sky130A
magscale 1 2
timestamp 1709454227
<< nwell >>
rect 4930 1030 5176 1088
rect 4930 1022 6004 1030
rect 8958 1022 9276 1092
rect 4930 1018 5176 1022
rect 8958 -638 9028 1022
rect 8958 -708 9208 -638
rect 11804 -706 11892 -638
<< pwell >>
rect 6428 -1096 6684 -1026
rect 8958 -1084 9158 -1026
rect 11800 -1084 11896 -1026
rect 6428 -1828 6504 -1096
rect 8958 -1754 9028 -1084
rect 8958 -1808 9268 -1754
<< locali >>
rect 6004 172 6152 228
rect 8514 132 8662 212
rect 11980 130 12136 220
rect 6116 -1898 6514 -1860
rect 8628 -1900 9028 -1854
rect 4118 -2590 4278 -2546
rect 3976 -2812 4154 -2778
<< viali >>
rect 5196 3376 5230 3422
rect 5196 3146 5230 3212
rect 8532 3148 8566 3228
rect 3834 2812 3872 2846
rect 4544 2526 4578 2596
rect 5482 1138 5548 1172
rect 8404 1140 8474 1174
rect 11514 1140 11580 1174
rect 6108 -2620 6156 -2568
rect 8626 -2626 8666 -2572
rect 12102 -2614 12140 -2554
rect 3942 -2812 3976 -2778
<< metal1 >>
rect 3798 3422 3998 3512
rect 5190 3422 5236 3434
rect 3798 3376 5196 3422
rect 5230 3376 5236 3422
rect 8764 3398 11534 3404
rect 8414 3396 11534 3398
rect 6622 3394 11534 3396
rect 3798 3312 3998 3376
rect 5190 3364 5236 3376
rect 5434 3332 11534 3394
rect 5434 3330 6278 3332
rect 3834 2852 3872 3312
rect 5190 3212 5236 3224
rect 5190 3208 5196 3212
rect 5230 3208 5236 3212
rect 5170 3152 5180 3208
rect 5248 3152 5258 3208
rect 5190 3146 5196 3152
rect 5230 3146 5236 3152
rect 5190 3134 5236 3146
rect 5380 3102 5390 3280
rect 5454 3102 5464 3280
rect 5574 3104 5584 3282
rect 5648 3104 5658 3282
rect 5766 3104 5776 3282
rect 5840 3104 5850 3282
rect 5958 3106 5968 3284
rect 6032 3106 6042 3284
rect 6148 3104 6158 3282
rect 6222 3104 6232 3282
rect 3822 2846 3884 2852
rect 3822 2812 3834 2846
rect 3872 2812 3884 2846
rect 3822 2806 3884 2812
rect 4266 2760 4772 2762
rect 4076 2692 4772 2760
rect 4022 2474 4032 2652
rect 4096 2474 4106 2652
rect 4214 2474 4224 2652
rect 4288 2474 4298 2652
rect 4406 2476 4416 2654
rect 4474 2588 4484 2654
rect 4538 2596 4584 2608
rect 4538 2588 4544 2596
rect 4474 2534 4544 2588
rect 4474 2476 4484 2534
rect 4538 2526 4544 2534
rect 4578 2526 4584 2596
rect 4538 2514 4584 2526
rect 4694 1662 4774 2692
rect 5284 1702 5294 1880
rect 5358 1702 5368 1880
rect 5478 1706 5488 1884
rect 5552 1706 5562 1884
rect 5668 1706 5678 1884
rect 5742 1706 5752 1884
rect 5858 1706 5868 1884
rect 5932 1706 5942 1884
rect 6050 1706 6060 1884
rect 6124 1706 6134 1884
rect 6242 1704 6252 1882
rect 6316 1704 6326 1882
rect 5294 1696 5354 1702
rect 4694 1650 6174 1662
rect 6372 1650 6418 3332
rect 6622 3328 8788 3332
rect 8414 3326 8788 3328
rect 6568 3104 6578 3282
rect 6642 3104 6652 3282
rect 6760 3102 6770 3280
rect 6834 3102 6844 3280
rect 6952 3104 6962 3282
rect 7026 3104 7036 3282
rect 7146 3104 7156 3282
rect 7220 3104 7230 3282
rect 7338 3104 7348 3282
rect 7412 3104 7422 3282
rect 7528 3102 7538 3280
rect 7602 3102 7612 3280
rect 7720 3104 7730 3282
rect 7794 3104 7804 3282
rect 7914 3104 7924 3282
rect 7988 3104 7998 3282
rect 8104 3104 8114 3282
rect 8178 3104 8188 3282
rect 8296 3104 8306 3282
rect 8370 3104 8380 3282
rect 8526 3228 8572 3240
rect 8526 3220 8532 3228
rect 8566 3220 8572 3228
rect 8506 3156 8516 3220
rect 8584 3156 8594 3220
rect 8526 3148 8532 3156
rect 8566 3148 8572 3156
rect 8526 3136 8572 3148
rect 8716 3106 8726 3284
rect 8790 3106 8800 3284
rect 8908 3102 8918 3280
rect 8982 3102 8992 3280
rect 9102 3104 9112 3282
rect 9176 3104 9186 3282
rect 9292 3104 9302 3282
rect 9366 3104 9376 3282
rect 9484 3104 9494 3282
rect 9558 3104 9568 3282
rect 9674 3104 9684 3282
rect 9748 3104 9758 3282
rect 9870 3102 9880 3280
rect 9944 3102 9954 3280
rect 10062 3104 10072 3282
rect 10136 3104 10146 3282
rect 10254 3104 10264 3282
rect 10328 3104 10338 3282
rect 10446 3102 10456 3280
rect 10520 3102 10530 3280
rect 10638 3104 10648 3282
rect 10712 3104 10722 3282
rect 10830 3104 10840 3282
rect 10904 3104 10914 3282
rect 11020 3104 11030 3282
rect 11094 3104 11104 3282
rect 11214 3104 11224 3282
rect 11288 3104 11298 3282
rect 11404 3104 11414 3282
rect 11478 3104 11488 3282
rect 6472 1704 6482 1882
rect 6546 1704 6556 1882
rect 6664 1704 6674 1882
rect 6738 1704 6748 1882
rect 6854 1704 6864 1882
rect 6928 1704 6938 1882
rect 7050 1704 7060 1882
rect 7124 1704 7134 1882
rect 7244 1706 7254 1884
rect 7318 1706 7328 1884
rect 7434 1704 7444 1882
rect 7508 1704 7518 1882
rect 7626 1704 7636 1882
rect 7700 1704 7710 1882
rect 7814 1704 7824 1882
rect 7888 1704 7898 1882
rect 8006 1706 8016 1884
rect 8080 1706 8090 1884
rect 8198 1704 8208 1882
rect 8272 1704 8282 1882
rect 8394 1702 8404 1880
rect 8468 1702 8478 1880
rect 8620 1704 8630 1882
rect 8694 1704 8704 1882
rect 8812 1702 8822 1880
rect 8886 1702 8896 1880
rect 9002 1704 9012 1882
rect 9076 1704 9086 1882
rect 9196 1704 9206 1882
rect 9270 1704 9280 1882
rect 9386 1702 9396 1880
rect 9460 1702 9470 1880
rect 9582 1704 9592 1882
rect 9656 1704 9666 1882
rect 9770 1706 9780 1884
rect 9844 1706 9854 1884
rect 9966 1706 9976 1884
rect 10040 1706 10050 1884
rect 10156 1704 10166 1882
rect 10230 1704 10240 1882
rect 10348 1704 10358 1882
rect 10422 1704 10432 1882
rect 10542 1704 10552 1882
rect 10616 1704 10626 1882
rect 10734 1702 10744 1888
rect 10808 1702 10818 1888
rect 10924 1704 10934 1890
rect 10998 1704 11008 1890
rect 11116 1706 11126 1892
rect 11190 1706 11200 1892
rect 11308 1706 11318 1892
rect 11382 1706 11392 1892
rect 11502 1704 11512 1890
rect 11576 1704 11586 1890
rect 6524 1652 8330 1658
rect 8670 1652 11440 1654
rect 6524 1650 11440 1652
rect 4694 1598 11440 1650
rect 4694 1584 5390 1598
rect 6524 1584 11440 1598
rect 3928 -926 3938 -820
rect 3996 -926 4006 -820
rect 4126 -926 4136 -820
rect 4194 -926 4204 -820
rect 4312 -926 4322 -820
rect 4380 -926 4390 -820
rect 4326 -976 4380 -926
rect 4694 -976 4774 1584
rect 8290 1582 11440 1584
rect 5472 1178 5482 1184
rect 5470 1132 5482 1178
rect 5548 1178 5558 1184
rect 5472 1128 5482 1132
rect 5548 1132 5560 1178
rect 5548 1128 5558 1132
rect 8390 1128 8400 1196
rect 8470 1180 8480 1196
rect 11514 1180 11580 1704
rect 8470 1174 8486 1180
rect 8474 1140 8486 1174
rect 8470 1134 8486 1140
rect 11502 1174 11592 1180
rect 11502 1140 11514 1174
rect 11580 1140 11592 1174
rect 11502 1134 11592 1140
rect 8470 1128 8480 1134
rect 4932 1086 6006 1088
rect 4890 1022 6006 1086
rect 6442 1022 8516 1092
rect 4890 1018 5178 1022
rect 4890 -642 4968 1018
rect 5022 872 5032 978
rect 5090 872 5100 978
rect 5214 872 5224 978
rect 5282 872 5292 978
rect 5408 872 5418 978
rect 5476 872 5486 978
rect 5598 872 5608 978
rect 5666 872 5676 978
rect 5790 870 5800 976
rect 5858 870 5868 976
rect 5982 872 5992 978
rect 6050 872 6060 978
rect 5118 -600 5128 -494
rect 5186 -600 5196 -494
rect 5310 -600 5320 -494
rect 5378 -600 5388 -494
rect 5502 -600 5512 -494
rect 5570 -600 5580 -494
rect 5694 -600 5704 -494
rect 5762 -600 5772 -494
rect 5886 -600 5896 -494
rect 5954 -600 5964 -494
rect 6444 -496 6512 1022
rect 6718 1020 8516 1022
rect 8958 1022 11992 1092
rect 6572 874 6582 980
rect 6640 874 6650 980
rect 6764 874 6774 980
rect 6832 874 6842 980
rect 6956 874 6966 980
rect 7024 874 7034 980
rect 7148 874 7158 980
rect 7216 874 7226 980
rect 7340 874 7350 980
rect 7408 874 7418 980
rect 7532 874 7542 980
rect 7600 874 7610 980
rect 7724 874 7734 980
rect 7792 874 7802 980
rect 7916 874 7926 980
rect 7984 874 7994 980
rect 8108 874 8118 980
rect 8176 874 8186 980
rect 8300 874 8310 980
rect 8368 874 8378 980
rect 8492 874 8502 980
rect 8560 874 8570 980
rect 8958 -490 9028 1022
rect 9086 874 9096 980
rect 9154 874 9164 980
rect 9278 874 9288 980
rect 9346 874 9356 980
rect 9470 872 9480 978
rect 9538 872 9548 978
rect 9662 872 9672 978
rect 9730 872 9740 978
rect 9852 874 9862 980
rect 9920 874 9930 980
rect 10046 874 10056 980
rect 10114 874 10124 980
rect 10238 874 10248 980
rect 10306 874 10316 980
rect 10430 874 10440 980
rect 10498 874 10508 980
rect 10622 874 10632 980
rect 10690 874 10700 980
rect 10814 874 10824 980
rect 10882 874 10892 980
rect 11006 874 11016 980
rect 11074 874 11084 980
rect 11200 874 11210 980
rect 11268 874 11278 980
rect 11390 874 11400 980
rect 11458 874 11468 980
rect 11582 874 11592 980
rect 11650 874 11660 980
rect 11774 876 11784 982
rect 11842 876 11852 982
rect 11966 874 11976 980
rect 12034 874 12044 980
rect 6430 -600 6440 -496
rect 6512 -600 6522 -496
rect 6670 -598 6680 -494
rect 6734 -598 6744 -494
rect 6862 -598 6872 -494
rect 6926 -598 6936 -494
rect 7054 -598 7064 -494
rect 7118 -598 7128 -494
rect 7246 -598 7256 -494
rect 7310 -598 7320 -494
rect 7438 -598 7448 -494
rect 7502 -598 7512 -494
rect 7630 -598 7640 -494
rect 7694 -598 7704 -494
rect 7822 -598 7832 -494
rect 7886 -598 7896 -494
rect 8014 -596 8024 -492
rect 8078 -596 8088 -492
rect 8206 -598 8216 -494
rect 8270 -598 8280 -494
rect 8398 -598 8408 -494
rect 8462 -598 8472 -494
rect 8950 -598 8960 -490
rect 9026 -598 9036 -490
rect 9182 -598 9192 -492
rect 9250 -598 9260 -492
rect 9374 -598 9384 -492
rect 9442 -598 9452 -492
rect 9566 -598 9576 -492
rect 9634 -598 9644 -492
rect 9756 -596 9766 -490
rect 9824 -596 9834 -490
rect 9950 -596 9960 -490
rect 10018 -596 10028 -490
rect 10142 -596 10152 -490
rect 10210 -596 10220 -490
rect 10334 -598 10344 -492
rect 10402 -598 10412 -492
rect 10524 -598 10534 -492
rect 10592 -598 10602 -492
rect 10716 -598 10726 -492
rect 10784 -598 10794 -492
rect 10908 -598 10918 -492
rect 10976 -598 10986 -492
rect 11102 -596 11112 -490
rect 11170 -596 11180 -490
rect 11294 -598 11304 -492
rect 11362 -598 11372 -492
rect 11486 -596 11496 -490
rect 11554 -596 11564 -490
rect 11678 -598 11688 -492
rect 11746 -598 11756 -492
rect 11870 -596 11880 -490
rect 11938 -596 11948 -490
rect 6444 -638 6512 -600
rect 8958 -638 9028 -598
rect 4890 -644 5146 -642
rect 5844 -644 5924 -640
rect 4890 -710 5924 -644
rect 6444 -708 8420 -638
rect 8958 -706 11892 -638
rect 8958 -708 11828 -706
rect 6444 -710 6696 -708
rect 5074 -712 5924 -710
rect 5844 -832 5924 -712
rect 5842 -834 5930 -832
rect 5842 -894 5852 -834
rect 5920 -894 5930 -834
rect 4310 -978 4774 -976
rect 3976 -1040 4774 -978
rect 3976 -1042 4432 -1040
rect 3796 -1340 3996 -1276
rect 3796 -1402 4620 -1340
rect 3796 -1476 3996 -1402
rect 3828 -2778 4028 -2644
rect 4080 -2674 4150 -1402
rect 4712 -1450 4774 -1040
rect 4310 -1566 4320 -1450
rect 4372 -1566 4382 -1450
rect 4502 -1566 4512 -1450
rect 4564 -1566 4574 -1450
rect 4698 -1566 4708 -1450
rect 4760 -1488 4774 -1450
rect 4890 -1022 5744 -1020
rect 5844 -1022 5924 -894
rect 4890 -1090 5924 -1022
rect 8346 -1026 8418 -708
rect 8958 -1026 9024 -708
rect 11970 -812 12170 -748
rect 11970 -890 12030 -812
rect 12112 -890 12170 -812
rect 11970 -948 12170 -890
rect 4760 -1566 4770 -1488
rect 4890 -1752 4962 -1090
rect 5054 -1092 5908 -1090
rect 5848 -1094 5908 -1092
rect 6438 -1096 8420 -1026
rect 8958 -1084 11896 -1026
rect 6438 -1130 6514 -1096
rect 5022 -1250 5032 -1134
rect 5084 -1250 5094 -1134
rect 5214 -1252 5224 -1136
rect 5276 -1252 5286 -1136
rect 5406 -1252 5416 -1136
rect 5468 -1252 5478 -1136
rect 5598 -1252 5608 -1136
rect 5660 -1252 5670 -1136
rect 5790 -1252 5800 -1136
rect 5852 -1252 5862 -1136
rect 5984 -1252 5994 -1136
rect 6046 -1252 6056 -1136
rect 6428 -1250 6438 -1130
rect 6522 -1250 6532 -1130
rect 5118 -1712 5128 -1596
rect 5180 -1712 5190 -1596
rect 5310 -1712 5320 -1596
rect 5372 -1712 5382 -1596
rect 5502 -1712 5512 -1596
rect 5564 -1712 5574 -1596
rect 5696 -1714 5706 -1598
rect 5758 -1714 5768 -1598
rect 5888 -1712 5898 -1596
rect 5950 -1712 5960 -1596
rect 4884 -1812 6004 -1752
rect 6438 -1760 6514 -1250
rect 6574 -1254 6584 -1138
rect 6636 -1254 6646 -1138
rect 6766 -1254 6776 -1138
rect 6828 -1254 6838 -1138
rect 6958 -1252 6968 -1136
rect 7020 -1252 7030 -1136
rect 7148 -1254 7158 -1138
rect 7210 -1254 7220 -1138
rect 7342 -1252 7352 -1136
rect 7404 -1252 7414 -1136
rect 7534 -1254 7544 -1138
rect 7596 -1254 7606 -1138
rect 7726 -1254 7736 -1138
rect 7788 -1254 7798 -1138
rect 7918 -1254 7928 -1138
rect 7980 -1254 7990 -1138
rect 8110 -1252 8120 -1136
rect 8172 -1252 8182 -1136
rect 8302 -1252 8312 -1136
rect 8364 -1252 8374 -1136
rect 8494 -1254 8504 -1138
rect 8556 -1254 8566 -1138
rect 8958 -1140 9028 -1084
rect 8954 -1250 8964 -1140
rect 9022 -1250 9032 -1140
rect 9086 -1234 9096 -1128
rect 9154 -1234 9164 -1128
rect 9278 -1232 9288 -1126
rect 9346 -1232 9356 -1126
rect 9470 -1232 9480 -1126
rect 9538 -1232 9548 -1126
rect 9662 -1234 9672 -1128
rect 9730 -1234 9740 -1128
rect 9852 -1234 9862 -1128
rect 9920 -1234 9930 -1128
rect 10046 -1234 10056 -1128
rect 10114 -1234 10124 -1128
rect 10236 -1234 10246 -1128
rect 10304 -1234 10314 -1128
rect 10428 -1232 10438 -1126
rect 10496 -1232 10506 -1126
rect 10622 -1234 10632 -1128
rect 10690 -1234 10700 -1128
rect 10814 -1232 10824 -1126
rect 10882 -1232 10892 -1126
rect 11004 -1234 11014 -1128
rect 11072 -1234 11082 -1128
rect 11198 -1232 11208 -1126
rect 11266 -1232 11276 -1126
rect 11392 -1234 11402 -1128
rect 11460 -1234 11470 -1128
rect 11582 -1232 11592 -1126
rect 11650 -1232 11660 -1126
rect 11776 -1234 11786 -1128
rect 11844 -1234 11854 -1128
rect 11966 -1234 11976 -1128
rect 12034 -1234 12044 -1128
rect 6670 -1716 6680 -1600
rect 6732 -1716 6742 -1600
rect 6862 -1714 6872 -1598
rect 6924 -1714 6934 -1598
rect 7054 -1714 7064 -1598
rect 7116 -1714 7126 -1598
rect 7246 -1714 7256 -1598
rect 7308 -1714 7318 -1598
rect 7438 -1714 7448 -1598
rect 7500 -1714 7510 -1598
rect 7632 -1714 7642 -1598
rect 7694 -1714 7704 -1598
rect 7822 -1714 7832 -1598
rect 7884 -1714 7894 -1598
rect 8012 -1716 8022 -1600
rect 8074 -1716 8084 -1600
rect 8208 -1712 8218 -1596
rect 8270 -1712 8280 -1596
rect 8396 -1712 8406 -1596
rect 8458 -1712 8468 -1596
rect 8958 -1754 9028 -1250
rect 9182 -1704 9192 -1598
rect 9250 -1704 9260 -1598
rect 9374 -1706 9384 -1600
rect 9442 -1706 9452 -1600
rect 9564 -1704 9574 -1598
rect 9632 -1704 9642 -1598
rect 9756 -1704 9766 -1598
rect 9824 -1704 9834 -1598
rect 9952 -1706 9962 -1600
rect 10020 -1706 10030 -1600
rect 10140 -1704 10150 -1598
rect 10208 -1704 10218 -1598
rect 10334 -1704 10344 -1598
rect 10402 -1704 10412 -1598
rect 10524 -1704 10534 -1598
rect 10592 -1704 10602 -1598
rect 10716 -1704 10726 -1598
rect 10784 -1704 10794 -1598
rect 10908 -1704 10918 -1598
rect 10976 -1704 10986 -1598
rect 11098 -1704 11108 -1598
rect 11166 -1704 11176 -1598
rect 11294 -1706 11304 -1600
rect 11362 -1706 11372 -1600
rect 11486 -1706 11496 -1600
rect 11554 -1706 11564 -1600
rect 11678 -1702 11688 -1596
rect 11746 -1702 11756 -1596
rect 11870 -1706 11880 -1600
rect 11938 -1706 11948 -1600
rect 9230 -1754 11994 -1752
rect 6720 -1760 8516 -1758
rect 6438 -1828 8516 -1760
rect 8958 -1808 11994 -1754
rect 5170 -1948 6006 -1940
rect 5170 -1952 8514 -1948
rect 9230 -1952 11992 -1934
rect 5170 -1996 11992 -1952
rect 5170 -2000 9294 -1996
rect 5170 -2004 8514 -2000
rect 5024 -2164 5034 -2048
rect 5086 -2164 5096 -2048
rect 5216 -2166 5226 -2050
rect 5278 -2166 5288 -2050
rect 5408 -2164 5418 -2048
rect 5470 -2164 5480 -2048
rect 5596 -2166 5606 -2050
rect 5658 -2166 5668 -2050
rect 5790 -2166 5800 -2050
rect 5852 -2166 5862 -2050
rect 5982 -2166 5992 -2050
rect 6044 -2166 6054 -2050
rect 4216 -2626 4226 -2510
rect 4278 -2626 4288 -2510
rect 4406 -2626 4416 -2510
rect 4468 -2626 4478 -2510
rect 4598 -2628 4608 -2512
rect 4660 -2628 4670 -2512
rect 5118 -2626 5128 -2510
rect 5180 -2626 5190 -2510
rect 5310 -2626 5320 -2510
rect 5372 -2626 5382 -2510
rect 5504 -2628 5514 -2512
rect 5566 -2628 5576 -2512
rect 5692 -2626 5702 -2510
rect 5754 -2626 5764 -2510
rect 5888 -2626 5898 -2510
rect 5950 -2626 5960 -2510
rect 6102 -2566 6162 -2556
rect 6084 -2620 6094 -2566
rect 6164 -2620 6174 -2566
rect 6102 -2632 6162 -2620
rect 4262 -2674 5098 -2672
rect 4080 -2680 5922 -2674
rect 6268 -2680 6360 -2004
rect 6722 -2008 8514 -2004
rect 6574 -2166 6584 -2050
rect 6636 -2166 6646 -2050
rect 6766 -2166 6776 -2050
rect 6828 -2166 6838 -2050
rect 6960 -2166 6970 -2050
rect 7022 -2166 7032 -2050
rect 7152 -2168 7162 -2052
rect 7214 -2168 7224 -2052
rect 7344 -2166 7354 -2050
rect 7406 -2166 7416 -2050
rect 7536 -2166 7546 -2050
rect 7598 -2166 7608 -2050
rect 7726 -2168 7736 -2052
rect 7788 -2168 7798 -2052
rect 7918 -2166 7928 -2050
rect 7980 -2166 7990 -2050
rect 8110 -2166 8120 -2050
rect 8172 -2166 8182 -2050
rect 8302 -2166 8312 -2050
rect 8364 -2166 8374 -2050
rect 8496 -2166 8506 -2050
rect 8558 -2166 8568 -2050
rect 9090 -2156 9100 -2040
rect 9152 -2156 9162 -2040
rect 9278 -2158 9288 -2042
rect 9340 -2158 9350 -2042
rect 9474 -2158 9484 -2042
rect 9536 -2158 9546 -2042
rect 9664 -2156 9674 -2040
rect 9726 -2156 9736 -2040
rect 9858 -2156 9868 -2040
rect 9920 -2156 9930 -2040
rect 10048 -2158 10058 -2042
rect 10110 -2158 10120 -2042
rect 10238 -2158 10248 -2042
rect 10300 -2158 10310 -2042
rect 10432 -2156 10442 -2040
rect 10494 -2156 10504 -2040
rect 10622 -2158 10632 -2042
rect 10684 -2158 10694 -2042
rect 10816 -2156 10826 -2040
rect 10878 -2156 10888 -2040
rect 11010 -2156 11020 -2040
rect 11072 -2156 11082 -2040
rect 11200 -2156 11210 -2040
rect 11262 -2156 11272 -2040
rect 11394 -2156 11404 -2040
rect 11456 -2156 11466 -2040
rect 11582 -2158 11592 -2042
rect 11644 -2158 11654 -2042
rect 11776 -2158 11786 -2042
rect 11838 -2158 11848 -2042
rect 11968 -2154 11978 -2038
rect 12030 -2154 12040 -2038
rect 6670 -2628 6680 -2512
rect 6732 -2628 6742 -2512
rect 6864 -2628 6874 -2512
rect 6926 -2628 6936 -2512
rect 7056 -2628 7066 -2512
rect 7118 -2628 7128 -2512
rect 7246 -2628 7256 -2512
rect 7308 -2628 7318 -2512
rect 7438 -2628 7448 -2512
rect 7500 -2628 7510 -2512
rect 7630 -2630 7640 -2514
rect 7692 -2630 7702 -2514
rect 7824 -2628 7834 -2512
rect 7886 -2628 7896 -2512
rect 8014 -2628 8024 -2512
rect 8076 -2628 8086 -2512
rect 8206 -2626 8216 -2510
rect 8268 -2626 8278 -2510
rect 8398 -2630 8408 -2514
rect 8460 -2630 8470 -2514
rect 8620 -2572 8672 -2560
rect 8604 -2626 8614 -2572
rect 8678 -2626 8688 -2572
rect 9184 -2618 9194 -2502
rect 9246 -2618 9256 -2502
rect 9376 -2618 9386 -2502
rect 9438 -2618 9448 -2502
rect 9568 -2620 9578 -2504
rect 9630 -2620 9640 -2504
rect 9762 -2618 9772 -2502
rect 9824 -2618 9834 -2502
rect 9950 -2620 9960 -2504
rect 10012 -2620 10022 -2504
rect 10144 -2620 10154 -2504
rect 10206 -2620 10216 -2504
rect 10334 -2620 10344 -2504
rect 10396 -2620 10406 -2504
rect 10528 -2620 10538 -2504
rect 10590 -2620 10600 -2504
rect 10720 -2620 10730 -2504
rect 10782 -2620 10792 -2504
rect 10914 -2618 10924 -2502
rect 10976 -2618 10986 -2502
rect 11102 -2620 11112 -2504
rect 11164 -2620 11174 -2504
rect 11296 -2618 11306 -2502
rect 11358 -2618 11368 -2502
rect 11488 -2620 11498 -2504
rect 11550 -2620 11560 -2504
rect 11678 -2618 11688 -2502
rect 11740 -2618 11750 -2502
rect 11874 -2620 11884 -2504
rect 11936 -2620 11946 -2504
rect 12096 -2554 12146 -2542
rect 12096 -2558 12102 -2554
rect 12140 -2558 12146 -2554
rect 12082 -2614 12092 -2558
rect 12148 -2614 12158 -2558
rect 12096 -2626 12146 -2614
rect 8620 -2638 8672 -2626
rect 9132 -2674 11894 -2660
rect 6620 -2680 11894 -2674
rect 4080 -2722 11894 -2680
rect 4080 -2730 9212 -2722
rect 4080 -2734 8424 -2730
rect 4262 -2736 8424 -2734
rect 5096 -2738 5922 -2736
rect 6620 -2750 8424 -2736
rect 3828 -2812 3942 -2778
rect 3976 -2812 4028 -2778
rect 3828 -2844 4028 -2812
<< via1 >>
rect 5180 3152 5196 3208
rect 5196 3152 5230 3208
rect 5230 3152 5248 3208
rect 5390 3102 5454 3280
rect 5584 3104 5648 3282
rect 5776 3104 5840 3282
rect 5968 3106 6032 3284
rect 6158 3104 6222 3282
rect 4032 2474 4096 2652
rect 4224 2474 4288 2652
rect 4416 2476 4474 2654
rect 5294 1702 5358 1880
rect 5488 1706 5552 1884
rect 5678 1706 5742 1884
rect 5868 1706 5932 1884
rect 6060 1706 6124 1884
rect 6252 1704 6316 1882
rect 6578 3104 6642 3282
rect 6770 3102 6834 3280
rect 6962 3104 7026 3282
rect 7156 3104 7220 3282
rect 7348 3104 7412 3282
rect 7538 3102 7602 3280
rect 7730 3104 7794 3282
rect 7924 3104 7988 3282
rect 8114 3104 8178 3282
rect 8306 3104 8370 3282
rect 8516 3156 8532 3220
rect 8532 3156 8566 3220
rect 8566 3156 8584 3220
rect 8726 3106 8790 3284
rect 8918 3102 8982 3280
rect 9112 3104 9176 3282
rect 9302 3104 9366 3282
rect 9494 3104 9558 3282
rect 9684 3104 9748 3282
rect 9880 3102 9944 3280
rect 10072 3104 10136 3282
rect 10264 3104 10328 3282
rect 10456 3102 10520 3280
rect 10648 3104 10712 3282
rect 10840 3104 10904 3282
rect 11030 3104 11094 3282
rect 11224 3104 11288 3282
rect 11414 3104 11478 3282
rect 6482 1704 6546 1882
rect 6674 1704 6738 1882
rect 6864 1704 6928 1882
rect 7060 1704 7124 1882
rect 7254 1706 7318 1884
rect 7444 1704 7508 1882
rect 7636 1704 7700 1882
rect 7824 1704 7888 1882
rect 8016 1706 8080 1884
rect 8208 1704 8272 1882
rect 8404 1702 8468 1880
rect 8630 1704 8694 1882
rect 8822 1702 8886 1880
rect 9012 1704 9076 1882
rect 9206 1704 9270 1882
rect 9396 1702 9460 1880
rect 9592 1704 9656 1882
rect 9780 1706 9844 1884
rect 9976 1706 10040 1884
rect 10166 1704 10230 1882
rect 10358 1704 10422 1882
rect 10552 1704 10616 1882
rect 10744 1702 10808 1888
rect 10934 1704 10998 1890
rect 11126 1706 11190 1892
rect 11318 1706 11382 1892
rect 11512 1704 11576 1890
rect 3938 -926 3996 -820
rect 4136 -926 4194 -820
rect 4322 -926 4380 -820
rect 5482 1172 5548 1184
rect 5482 1138 5548 1172
rect 5482 1128 5548 1138
rect 8400 1174 8470 1196
rect 8400 1140 8404 1174
rect 8404 1140 8470 1174
rect 8400 1128 8470 1140
rect 5032 872 5090 978
rect 5224 872 5282 978
rect 5418 872 5476 978
rect 5608 872 5666 978
rect 5800 870 5858 976
rect 5992 872 6050 978
rect 5128 -600 5186 -494
rect 5320 -600 5378 -494
rect 5512 -600 5570 -494
rect 5704 -600 5762 -494
rect 5896 -600 5954 -494
rect 6582 874 6640 980
rect 6774 874 6832 980
rect 6966 874 7024 980
rect 7158 874 7216 980
rect 7350 874 7408 980
rect 7542 874 7600 980
rect 7734 874 7792 980
rect 7926 874 7984 980
rect 8118 874 8176 980
rect 8310 874 8368 980
rect 8502 874 8560 980
rect 9096 874 9154 980
rect 9288 874 9346 980
rect 9480 872 9538 978
rect 9672 872 9730 978
rect 9862 874 9920 980
rect 10056 874 10114 980
rect 10248 874 10306 980
rect 10440 874 10498 980
rect 10632 874 10690 980
rect 10824 874 10882 980
rect 11016 874 11074 980
rect 11210 874 11268 980
rect 11400 874 11458 980
rect 11592 874 11650 980
rect 11784 876 11842 982
rect 11976 874 12034 980
rect 6440 -600 6512 -496
rect 6680 -598 6734 -494
rect 6872 -598 6926 -494
rect 7064 -598 7118 -494
rect 7256 -598 7310 -494
rect 7448 -598 7502 -494
rect 7640 -598 7694 -494
rect 7832 -598 7886 -494
rect 8024 -596 8078 -492
rect 8216 -598 8270 -494
rect 8408 -598 8462 -494
rect 8960 -598 9026 -490
rect 9192 -598 9250 -492
rect 9384 -598 9442 -492
rect 9576 -598 9634 -492
rect 9766 -596 9824 -490
rect 9960 -596 10018 -490
rect 10152 -596 10210 -490
rect 10344 -598 10402 -492
rect 10534 -598 10592 -492
rect 10726 -598 10784 -492
rect 10918 -598 10976 -492
rect 11112 -596 11170 -490
rect 11304 -598 11362 -492
rect 11496 -596 11554 -490
rect 11688 -598 11746 -492
rect 11880 -596 11938 -490
rect 5852 -894 5920 -834
rect 4320 -1566 4372 -1450
rect 4512 -1566 4564 -1450
rect 4708 -1566 4760 -1450
rect 12030 -890 12112 -812
rect 5032 -1250 5084 -1134
rect 5224 -1252 5276 -1136
rect 5416 -1252 5468 -1136
rect 5608 -1252 5660 -1136
rect 5800 -1252 5852 -1136
rect 5994 -1252 6046 -1136
rect 6438 -1250 6522 -1130
rect 5128 -1712 5180 -1596
rect 5320 -1712 5372 -1596
rect 5512 -1712 5564 -1596
rect 5706 -1714 5758 -1598
rect 5898 -1712 5950 -1596
rect 6584 -1254 6636 -1138
rect 6776 -1254 6828 -1138
rect 6968 -1252 7020 -1136
rect 7158 -1254 7210 -1138
rect 7352 -1252 7404 -1136
rect 7544 -1254 7596 -1138
rect 7736 -1254 7788 -1138
rect 7928 -1254 7980 -1138
rect 8120 -1252 8172 -1136
rect 8312 -1252 8364 -1136
rect 8504 -1254 8556 -1138
rect 8964 -1250 9022 -1140
rect 9096 -1234 9154 -1128
rect 9288 -1232 9346 -1126
rect 9480 -1232 9538 -1126
rect 9672 -1234 9730 -1128
rect 9862 -1234 9920 -1128
rect 10056 -1234 10114 -1128
rect 10246 -1234 10304 -1128
rect 10438 -1232 10496 -1126
rect 10632 -1234 10690 -1128
rect 10824 -1232 10882 -1126
rect 11014 -1234 11072 -1128
rect 11208 -1232 11266 -1126
rect 11402 -1234 11460 -1128
rect 11592 -1232 11650 -1126
rect 11786 -1234 11844 -1128
rect 11976 -1234 12034 -1128
rect 6680 -1716 6732 -1600
rect 6872 -1714 6924 -1598
rect 7064 -1714 7116 -1598
rect 7256 -1714 7308 -1598
rect 7448 -1714 7500 -1598
rect 7642 -1714 7694 -1598
rect 7832 -1714 7884 -1598
rect 8022 -1716 8074 -1600
rect 8218 -1712 8270 -1596
rect 8406 -1712 8458 -1596
rect 9192 -1704 9250 -1598
rect 9384 -1706 9442 -1600
rect 9574 -1704 9632 -1598
rect 9766 -1704 9824 -1598
rect 9962 -1706 10020 -1600
rect 10150 -1704 10208 -1598
rect 10344 -1704 10402 -1598
rect 10534 -1704 10592 -1598
rect 10726 -1704 10784 -1598
rect 10918 -1704 10976 -1598
rect 11108 -1704 11166 -1598
rect 11304 -1706 11362 -1600
rect 11496 -1706 11554 -1600
rect 11688 -1702 11746 -1596
rect 11880 -1706 11938 -1600
rect 5034 -2164 5086 -2048
rect 5226 -2166 5278 -2050
rect 5418 -2164 5470 -2048
rect 5606 -2166 5658 -2050
rect 5800 -2166 5852 -2050
rect 5992 -2166 6044 -2050
rect 4226 -2626 4278 -2510
rect 4416 -2626 4468 -2510
rect 4608 -2628 4660 -2512
rect 5128 -2626 5180 -2510
rect 5320 -2626 5372 -2510
rect 5514 -2628 5566 -2512
rect 5702 -2626 5754 -2510
rect 5898 -2626 5950 -2510
rect 6094 -2568 6164 -2566
rect 6094 -2620 6108 -2568
rect 6108 -2620 6156 -2568
rect 6156 -2620 6164 -2568
rect 6584 -2166 6636 -2050
rect 6776 -2166 6828 -2050
rect 6970 -2166 7022 -2050
rect 7162 -2168 7214 -2052
rect 7354 -2166 7406 -2050
rect 7546 -2166 7598 -2050
rect 7736 -2168 7788 -2052
rect 7928 -2166 7980 -2050
rect 8120 -2166 8172 -2050
rect 8312 -2166 8364 -2050
rect 8506 -2166 8558 -2050
rect 9100 -2156 9152 -2040
rect 9288 -2158 9340 -2042
rect 9484 -2158 9536 -2042
rect 9674 -2156 9726 -2040
rect 9868 -2156 9920 -2040
rect 10058 -2158 10110 -2042
rect 10248 -2158 10300 -2042
rect 10442 -2156 10494 -2040
rect 10632 -2158 10684 -2042
rect 10826 -2156 10878 -2040
rect 11020 -2156 11072 -2040
rect 11210 -2156 11262 -2040
rect 11404 -2156 11456 -2040
rect 11592 -2158 11644 -2042
rect 11786 -2158 11838 -2042
rect 11978 -2154 12030 -2038
rect 6680 -2628 6732 -2512
rect 6874 -2628 6926 -2512
rect 7066 -2628 7118 -2512
rect 7256 -2628 7308 -2512
rect 7448 -2628 7500 -2512
rect 7640 -2630 7692 -2514
rect 7834 -2628 7886 -2512
rect 8024 -2628 8076 -2512
rect 8216 -2626 8268 -2510
rect 8408 -2630 8460 -2514
rect 8614 -2626 8626 -2572
rect 8626 -2626 8666 -2572
rect 8666 -2626 8678 -2572
rect 9194 -2618 9246 -2502
rect 9386 -2618 9438 -2502
rect 9578 -2620 9630 -2504
rect 9772 -2618 9824 -2502
rect 9960 -2620 10012 -2504
rect 10154 -2620 10206 -2504
rect 10344 -2620 10396 -2504
rect 10538 -2620 10590 -2504
rect 10730 -2620 10782 -2504
rect 10924 -2618 10976 -2502
rect 11112 -2620 11164 -2504
rect 11306 -2618 11358 -2502
rect 11498 -2620 11550 -2504
rect 11688 -2618 11740 -2502
rect 11884 -2620 11936 -2504
rect 12092 -2614 12102 -2558
rect 12102 -2614 12140 -2558
rect 12140 -2614 12148 -2558
<< metal2 >>
rect 5390 3284 5454 3290
rect 5584 3284 5648 3292
rect 5776 3284 5840 3292
rect 5968 3284 6032 3294
rect 6158 3284 6222 3292
rect 5382 3282 5968 3284
rect 5382 3280 5584 3282
rect 5180 3208 5248 3218
rect 5382 3208 5390 3280
rect 5248 3152 5390 3208
rect 5180 3142 5248 3152
rect 5382 3102 5390 3152
rect 5454 3104 5584 3280
rect 5648 3104 5776 3282
rect 5840 3106 5968 3282
rect 6032 3282 6230 3284
rect 6032 3106 6158 3282
rect 5840 3104 6158 3106
rect 6222 3104 6230 3282
rect 5454 3102 6230 3104
rect 5382 3098 6230 3102
rect 6564 3282 8382 3296
rect 6564 3104 6578 3282
rect 6642 3280 6962 3282
rect 6642 3104 6770 3280
rect 6564 3102 6770 3104
rect 6834 3104 6962 3280
rect 7026 3104 7156 3282
rect 7220 3104 7348 3282
rect 7412 3280 7730 3282
rect 7412 3104 7538 3280
rect 6834 3102 7538 3104
rect 7602 3104 7730 3280
rect 7794 3104 7924 3282
rect 7988 3104 8114 3282
rect 8178 3104 8306 3282
rect 8370 3220 8382 3282
rect 8712 3284 11490 3298
rect 8516 3220 8584 3230
rect 8712 3220 8726 3284
rect 8370 3156 8516 3220
rect 8584 3156 8726 3220
rect 8370 3104 8382 3156
rect 8516 3146 8584 3156
rect 7602 3102 8382 3104
rect 5390 3092 5454 3098
rect 5584 3094 5648 3098
rect 5776 3094 5840 3098
rect 5968 3096 6032 3098
rect 6158 3094 6222 3098
rect 6564 3092 8382 3102
rect 8712 3106 8726 3156
rect 8790 3282 11490 3284
rect 8790 3280 9112 3282
rect 8790 3106 8918 3280
rect 8712 3102 8918 3106
rect 8982 3104 9112 3280
rect 9176 3104 9302 3282
rect 9366 3104 9494 3282
rect 9558 3104 9684 3282
rect 9748 3280 10072 3282
rect 9748 3104 9880 3280
rect 8982 3102 9880 3104
rect 9944 3104 10072 3280
rect 10136 3104 10264 3282
rect 10328 3280 10648 3282
rect 10328 3104 10456 3280
rect 9944 3102 10456 3104
rect 10520 3104 10648 3280
rect 10712 3104 10840 3282
rect 10904 3104 11030 3282
rect 11094 3104 11224 3282
rect 11288 3104 11414 3282
rect 11478 3104 11490 3282
rect 10520 3102 11490 3104
rect 8712 3100 11490 3102
rect 8726 3096 8790 3100
rect 8918 3092 8982 3100
rect 9112 3094 9176 3100
rect 9302 3094 9366 3100
rect 9494 3094 9558 3100
rect 9684 3094 9748 3100
rect 9880 3092 9944 3100
rect 10072 3094 10136 3100
rect 10264 3094 10328 3100
rect 10456 3092 10520 3100
rect 10648 3094 10712 3100
rect 10840 3094 10904 3100
rect 11030 3094 11094 3100
rect 11224 3094 11288 3100
rect 11414 3094 11478 3100
rect 4416 2662 4474 2664
rect 4030 2654 4476 2662
rect 4030 2652 4416 2654
rect 4030 2474 4032 2652
rect 4096 2474 4224 2652
rect 4288 2476 4416 2652
rect 4474 2476 4476 2654
rect 4288 2474 4476 2476
rect 4030 2466 4476 2474
rect 4032 2464 4096 2466
rect 4224 2464 4288 2466
rect 10744 1896 10808 1898
rect 10934 1896 10998 1900
rect 11126 1896 11190 1902
rect 11318 1896 11382 1902
rect 11512 1896 11576 1900
rect 5294 1882 5358 1890
rect 5488 1884 5552 1894
rect 5294 1880 5488 1882
rect 5358 1706 5488 1880
rect 5678 1884 5742 1894
rect 5552 1706 5678 1882
rect 5868 1884 5932 1894
rect 5742 1706 5868 1882
rect 6060 1884 6124 1894
rect 5932 1706 6060 1882
rect 6252 1882 6316 1892
rect 6482 1886 6546 1892
rect 6674 1886 6738 1892
rect 6864 1886 6928 1892
rect 7060 1886 7124 1892
rect 7254 1886 7318 1894
rect 7444 1886 7508 1892
rect 7636 1886 7700 1892
rect 7824 1886 7888 1892
rect 8016 1886 8080 1894
rect 8616 1892 11588 1896
rect 8208 1886 8272 1892
rect 8616 1890 11126 1892
rect 8404 1886 8468 1890
rect 8616 1888 10934 1890
rect 6472 1884 8472 1886
rect 6472 1882 7254 1884
rect 6124 1706 6252 1882
rect 5358 1704 6252 1706
rect 6316 1704 6322 1882
rect 5358 1702 6322 1704
rect 5294 1698 6322 1702
rect 6472 1704 6482 1882
rect 6546 1704 6674 1882
rect 6738 1704 6864 1882
rect 6928 1704 7060 1882
rect 7124 1706 7254 1882
rect 7318 1882 8016 1884
rect 7318 1706 7444 1882
rect 7124 1704 7444 1706
rect 7508 1704 7636 1882
rect 7700 1704 7824 1882
rect 7888 1706 8016 1882
rect 8080 1882 8472 1884
rect 8080 1706 8208 1882
rect 7888 1704 8208 1706
rect 8272 1880 8472 1882
rect 8272 1704 8404 1880
rect 6472 1702 8404 1704
rect 8468 1702 8472 1880
rect 5294 1692 5358 1698
rect 5482 1696 5552 1698
rect 5678 1696 5742 1698
rect 5868 1696 5932 1698
rect 6060 1696 6124 1698
rect 5482 1194 5546 1696
rect 6252 1694 6316 1698
rect 6472 1696 8472 1702
rect 8616 1884 10744 1888
rect 8616 1882 9780 1884
rect 8616 1704 8630 1882
rect 8694 1880 9012 1882
rect 8694 1704 8822 1880
rect 8616 1702 8822 1704
rect 8886 1704 9012 1880
rect 9076 1704 9206 1882
rect 9270 1880 9592 1882
rect 9270 1704 9396 1880
rect 8886 1702 9396 1704
rect 9460 1704 9592 1880
rect 9656 1706 9780 1882
rect 9844 1706 9976 1884
rect 10040 1882 10744 1884
rect 10040 1706 10166 1882
rect 9656 1704 10166 1706
rect 10230 1704 10358 1882
rect 10422 1704 10552 1882
rect 10616 1704 10744 1882
rect 9460 1702 10744 1704
rect 10808 1704 10934 1888
rect 10998 1706 11126 1890
rect 11190 1706 11318 1892
rect 11382 1890 11588 1892
rect 11382 1706 11512 1890
rect 10998 1704 11512 1706
rect 11576 1704 11588 1890
rect 10808 1702 11588 1704
rect 6482 1694 6546 1696
rect 6674 1694 6738 1696
rect 6864 1694 6928 1696
rect 7060 1694 7124 1696
rect 7444 1694 7508 1696
rect 7636 1694 7700 1696
rect 7824 1694 7888 1696
rect 8208 1694 8272 1696
rect 8400 1692 8468 1696
rect 8616 1694 11588 1702
rect 8822 1692 8886 1694
rect 9396 1692 9460 1694
rect 10744 1692 10808 1694
rect 8400 1206 8464 1692
rect 8400 1196 8470 1206
rect 5482 1184 5548 1194
rect 5482 1118 5548 1128
rect 8400 1118 8470 1128
rect 5022 978 6060 990
rect 5022 872 5032 978
rect 5090 872 5224 978
rect 5282 872 5418 978
rect 5476 872 5608 978
rect 5666 976 5992 978
rect 5666 872 5800 976
rect 5022 870 5800 872
rect 5858 872 5992 976
rect 6050 872 6060 978
rect 5858 870 6060 872
rect 5022 862 6060 870
rect 6566 980 8576 994
rect 9096 988 9154 990
rect 9288 988 9346 990
rect 9862 988 9920 990
rect 10056 988 10114 990
rect 10248 988 10306 990
rect 10440 988 10498 990
rect 10632 988 10690 990
rect 10824 988 10882 990
rect 11016 988 11074 990
rect 11210 988 11268 990
rect 11400 988 11458 990
rect 11592 988 11650 990
rect 11784 988 11842 992
rect 11976 988 12034 990
rect 6566 874 6582 980
rect 6640 874 6774 980
rect 6832 874 6966 980
rect 7024 874 7158 980
rect 7216 874 7350 980
rect 7408 874 7542 980
rect 7600 874 7734 980
rect 7792 874 7926 980
rect 7984 874 8118 980
rect 8176 874 8310 980
rect 8368 874 8502 980
rect 8560 874 8576 980
rect 9082 982 12046 988
rect 9082 980 11784 982
rect 9082 874 9096 980
rect 9154 874 9288 980
rect 9346 978 9862 980
rect 9346 874 9480 978
rect 6566 868 8576 874
rect 6582 864 6640 868
rect 6774 864 6832 868
rect 6966 864 7024 868
rect 7158 864 7216 868
rect 7350 864 7408 868
rect 7542 864 7600 868
rect 7734 864 7792 868
rect 7926 864 7984 868
rect 8118 864 8176 868
rect 8310 864 8368 868
rect 8502 864 8560 868
rect 9096 864 9154 874
rect 9288 864 9346 874
rect 9538 874 9672 978
rect 9480 862 9538 872
rect 9730 874 9862 978
rect 9920 874 10056 980
rect 10114 874 10248 980
rect 10306 874 10440 980
rect 10498 874 10632 980
rect 10690 874 10824 980
rect 10882 874 11016 980
rect 11074 874 11210 980
rect 11268 874 11400 980
rect 11458 874 11592 980
rect 11650 876 11784 980
rect 11842 980 12046 982
rect 11842 876 11976 980
rect 11650 874 11976 876
rect 12034 874 12046 980
rect 9672 862 9730 872
rect 9862 864 9920 874
rect 10056 864 10114 874
rect 10248 864 10306 874
rect 10440 864 10498 874
rect 10632 864 10690 874
rect 10824 864 10882 874
rect 11016 864 11074 874
rect 11210 864 11268 874
rect 11400 864 11458 874
rect 11592 864 11650 874
rect 11784 866 11842 874
rect 11976 864 12034 874
rect 5800 860 5858 862
rect 5128 -492 5186 -484
rect 5320 -492 5378 -484
rect 5512 -492 5570 -484
rect 5704 -492 5762 -484
rect 5896 -492 5954 -484
rect 5116 -494 5964 -492
rect 5116 -600 5128 -494
rect 5186 -600 5320 -494
rect 5378 -600 5512 -494
rect 5570 -600 5704 -494
rect 5762 -600 5896 -494
rect 5954 -498 5964 -494
rect 6440 -496 6512 -486
rect 5954 -600 6440 -498
rect 6666 -490 8468 -482
rect 8960 -490 9026 -480
rect 6666 -492 8960 -490
rect 6666 -494 8024 -492
rect 6512 -600 6514 -498
rect 6666 -596 6680 -494
rect 5128 -610 5186 -600
rect 5320 -610 5378 -600
rect 5512 -610 5570 -600
rect 5704 -610 5762 -600
rect 5896 -604 6514 -600
rect 6734 -596 6872 -494
rect 5896 -610 5954 -604
rect 6440 -610 6512 -604
rect 6680 -608 6734 -598
rect 6926 -596 7064 -494
rect 6872 -608 6926 -598
rect 7118 -596 7256 -494
rect 7064 -608 7118 -598
rect 7310 -596 7448 -494
rect 7256 -608 7310 -598
rect 7502 -596 7640 -494
rect 7448 -608 7502 -598
rect 7694 -596 7832 -494
rect 7640 -608 7694 -598
rect 7886 -596 8024 -494
rect 8078 -494 8960 -492
rect 8078 -596 8216 -494
rect 7832 -608 7886 -598
rect 8024 -606 8078 -596
rect 8270 -596 8408 -494
rect 8216 -608 8270 -598
rect 8462 -594 8960 -494
rect 8462 -596 8468 -594
rect 8408 -608 8462 -598
rect 8960 -608 9026 -598
rect 9182 -490 11942 -478
rect 9182 -492 9766 -490
rect 9182 -598 9192 -492
rect 9250 -598 9384 -492
rect 9442 -598 9576 -492
rect 9634 -596 9766 -492
rect 9824 -596 9960 -490
rect 10018 -596 10152 -490
rect 10210 -492 11112 -490
rect 10210 -596 10344 -492
rect 9634 -598 10344 -596
rect 10402 -598 10534 -492
rect 10592 -598 10726 -492
rect 10784 -598 10918 -492
rect 10976 -596 11112 -492
rect 11170 -492 11496 -490
rect 11170 -596 11304 -492
rect 10976 -598 11304 -596
rect 11362 -596 11496 -492
rect 11554 -492 11880 -490
rect 11554 -596 11688 -492
rect 11362 -598 11688 -596
rect 11746 -596 11880 -492
rect 11938 -534 11942 -490
rect 11938 -594 12116 -534
rect 11938 -596 11942 -594
rect 11746 -598 11942 -596
rect 9182 -604 11942 -598
rect 9192 -608 9250 -604
rect 9384 -608 9442 -604
rect 9576 -608 9634 -604
rect 9766 -606 9824 -604
rect 9960 -606 10018 -604
rect 10152 -606 10210 -604
rect 10344 -608 10402 -604
rect 10534 -608 10592 -604
rect 10726 -608 10784 -604
rect 10918 -608 10976 -604
rect 11112 -606 11170 -604
rect 11304 -608 11362 -604
rect 11496 -606 11554 -604
rect 11688 -608 11746 -604
rect 11880 -606 11938 -604
rect 12034 -800 12106 -594
rect 3938 -812 3996 -810
rect 4136 -812 4194 -810
rect 4322 -812 4380 -810
rect 12030 -812 12112 -800
rect 3936 -820 4386 -812
rect 3936 -926 3938 -820
rect 3996 -926 4136 -820
rect 4194 -926 4322 -820
rect 4380 -926 4386 -820
rect 5842 -834 12030 -820
rect 5842 -894 5852 -834
rect 5920 -890 12030 -834
rect 12112 -890 12116 -820
rect 5920 -894 12116 -890
rect 5842 -898 12116 -894
rect 5852 -904 5920 -898
rect 3936 -936 4386 -926
rect 5032 -1134 5084 -1124
rect 5026 -1250 5032 -1136
rect 5224 -1136 5276 -1126
rect 5416 -1136 5468 -1126
rect 5608 -1136 5660 -1126
rect 5800 -1136 5852 -1126
rect 5994 -1132 6046 -1126
rect 6438 -1130 6522 -1120
rect 9096 -1126 9154 -1118
rect 9288 -1126 9346 -1116
rect 9480 -1126 9538 -1116
rect 9672 -1126 9730 -1118
rect 9862 -1126 9920 -1118
rect 10056 -1126 10114 -1118
rect 10246 -1126 10304 -1118
rect 10438 -1126 10496 -1116
rect 10632 -1126 10690 -1118
rect 10824 -1126 10882 -1116
rect 11014 -1126 11072 -1118
rect 11208 -1126 11266 -1116
rect 11402 -1126 11460 -1118
rect 11592 -1126 11650 -1116
rect 12030 -1118 12112 -898
rect 11786 -1126 11844 -1118
rect 11976 -1126 12112 -1118
rect 5994 -1136 6438 -1132
rect 5084 -1250 5224 -1136
rect 5026 -1252 5224 -1250
rect 5276 -1252 5416 -1136
rect 5468 -1252 5608 -1136
rect 5660 -1252 5800 -1136
rect 5852 -1252 5994 -1136
rect 6046 -1250 6438 -1136
rect 6046 -1252 6522 -1250
rect 5032 -1260 5084 -1252
rect 5224 -1262 5276 -1252
rect 5416 -1262 5468 -1252
rect 5608 -1262 5660 -1252
rect 5800 -1262 5852 -1252
rect 5994 -1262 6046 -1252
rect 6438 -1260 6522 -1252
rect 6584 -1138 6636 -1128
rect 6776 -1138 6828 -1128
rect 6636 -1252 6776 -1140
rect 6584 -1264 6636 -1254
rect 6968 -1136 7020 -1126
rect 6828 -1252 6968 -1140
rect 7158 -1138 7210 -1128
rect 7020 -1252 7158 -1140
rect 6776 -1264 6828 -1254
rect 6968 -1262 7020 -1252
rect 7352 -1136 7404 -1126
rect 7210 -1252 7352 -1140
rect 7544 -1138 7596 -1128
rect 7404 -1252 7544 -1140
rect 7158 -1264 7210 -1254
rect 7352 -1262 7404 -1252
rect 7736 -1138 7788 -1128
rect 7596 -1252 7736 -1140
rect 7544 -1264 7596 -1254
rect 7928 -1138 7980 -1128
rect 7788 -1252 7928 -1140
rect 7736 -1264 7788 -1254
rect 8120 -1136 8172 -1126
rect 7980 -1252 8120 -1140
rect 8312 -1136 8364 -1126
rect 9080 -1128 9288 -1126
rect 8172 -1252 8312 -1140
rect 8504 -1130 8556 -1128
rect 8504 -1138 9026 -1130
rect 8364 -1252 8504 -1140
rect 7928 -1264 7980 -1254
rect 8120 -1262 8172 -1252
rect 8312 -1262 8364 -1252
rect 8556 -1140 9026 -1138
rect 8556 -1250 8964 -1140
rect 9022 -1250 9026 -1140
rect 9080 -1234 9096 -1128
rect 9154 -1232 9288 -1128
rect 9346 -1232 9480 -1126
rect 9538 -1128 10438 -1126
rect 9538 -1232 9672 -1128
rect 9154 -1234 9672 -1232
rect 9730 -1234 9862 -1128
rect 9920 -1234 10056 -1128
rect 10114 -1234 10246 -1128
rect 10304 -1232 10438 -1128
rect 10496 -1128 10824 -1126
rect 10496 -1232 10632 -1128
rect 10304 -1234 10632 -1232
rect 10690 -1232 10824 -1128
rect 10882 -1128 11208 -1126
rect 10882 -1232 11014 -1128
rect 10690 -1234 11014 -1232
rect 11072 -1232 11208 -1128
rect 11266 -1128 11592 -1126
rect 11266 -1232 11402 -1128
rect 11072 -1234 11402 -1232
rect 11460 -1232 11592 -1128
rect 11650 -1128 12112 -1126
rect 11650 -1232 11786 -1128
rect 11460 -1234 11786 -1232
rect 11844 -1234 11976 -1128
rect 12034 -1170 12112 -1128
rect 12034 -1234 12044 -1170
rect 9080 -1236 12044 -1234
rect 9096 -1244 9154 -1236
rect 9288 -1242 9346 -1236
rect 9480 -1242 9538 -1236
rect 9672 -1244 9730 -1236
rect 9862 -1244 9920 -1236
rect 10056 -1244 10114 -1236
rect 10246 -1244 10304 -1236
rect 10438 -1242 10496 -1236
rect 10632 -1244 10690 -1236
rect 10824 -1242 10882 -1236
rect 11014 -1244 11072 -1236
rect 11208 -1242 11266 -1236
rect 11402 -1244 11460 -1236
rect 11592 -1242 11650 -1236
rect 11786 -1244 11844 -1236
rect 11976 -1244 12034 -1236
rect 8556 -1252 9026 -1250
rect 8504 -1264 8556 -1254
rect 8964 -1260 9022 -1252
rect 4320 -1446 4372 -1440
rect 4512 -1446 4564 -1440
rect 4708 -1446 4760 -1440
rect 4312 -1450 4770 -1446
rect 4312 -1566 4320 -1450
rect 4372 -1566 4512 -1450
rect 4564 -1566 4708 -1450
rect 4760 -1566 4770 -1450
rect 4312 -1568 4770 -1566
rect 4320 -1576 4372 -1568
rect 4512 -1576 4564 -1568
rect 4708 -1576 4760 -1568
rect 5128 -1588 5180 -1586
rect 5320 -1588 5372 -1586
rect 5512 -1588 5564 -1586
rect 5898 -1588 5950 -1586
rect 5120 -1596 5954 -1588
rect 5120 -1710 5128 -1596
rect 5180 -1710 5320 -1596
rect 5128 -1722 5180 -1712
rect 5372 -1710 5512 -1596
rect 5320 -1722 5372 -1712
rect 5564 -1598 5898 -1596
rect 5564 -1710 5706 -1598
rect 5512 -1722 5564 -1712
rect 5758 -1710 5898 -1598
rect 5706 -1724 5758 -1714
rect 5876 -1712 5898 -1710
rect 5950 -1712 5954 -1596
rect 5034 -2048 5086 -2038
rect 5022 -2164 5034 -2050
rect 5226 -2050 5278 -2040
rect 5418 -2048 5470 -2038
rect 5876 -2040 5954 -1712
rect 6680 -1594 6732 -1590
rect 6872 -1594 6924 -1588
rect 7064 -1594 7116 -1588
rect 7256 -1594 7308 -1588
rect 7448 -1594 7500 -1588
rect 7642 -1594 7694 -1588
rect 7832 -1594 7884 -1588
rect 8022 -1594 8074 -1590
rect 8218 -1594 8270 -1586
rect 8406 -1594 8458 -1586
rect 6680 -1596 8458 -1594
rect 6680 -1598 8218 -1596
rect 6680 -1600 6872 -1598
rect 6732 -1714 6872 -1600
rect 6924 -1714 7064 -1598
rect 7116 -1714 7256 -1598
rect 7308 -1714 7448 -1598
rect 7500 -1714 7642 -1598
rect 7694 -1714 7832 -1598
rect 7884 -1600 8218 -1598
rect 7884 -1714 8022 -1600
rect 6732 -1716 8022 -1714
rect 8074 -1712 8218 -1600
rect 8270 -1712 8406 -1596
rect 9182 -1596 11940 -1586
rect 9182 -1598 11688 -1596
rect 9182 -1704 9192 -1598
rect 9250 -1600 9574 -1598
rect 9250 -1704 9384 -1600
rect 9182 -1706 9384 -1704
rect 9442 -1704 9574 -1600
rect 9632 -1704 9766 -1598
rect 9824 -1600 10150 -1598
rect 9824 -1704 9962 -1600
rect 9442 -1706 9962 -1704
rect 10020 -1704 10150 -1600
rect 10208 -1704 10344 -1598
rect 10402 -1704 10534 -1598
rect 10592 -1704 10726 -1598
rect 10784 -1704 10918 -1598
rect 10976 -1704 11108 -1598
rect 11166 -1600 11688 -1598
rect 11166 -1704 11304 -1600
rect 10020 -1706 11304 -1704
rect 11362 -1706 11496 -1600
rect 11554 -1702 11688 -1600
rect 11746 -1600 11940 -1596
rect 11746 -1702 11880 -1600
rect 11554 -1706 11880 -1702
rect 11938 -1706 11940 -1600
rect 9182 -1708 11940 -1706
rect 8074 -1716 8458 -1712
rect 9192 -1714 9250 -1708
rect 9384 -1716 9442 -1708
rect 9574 -1714 9632 -1708
rect 9766 -1714 9824 -1708
rect 9962 -1716 10020 -1708
rect 10150 -1714 10208 -1708
rect 10344 -1714 10402 -1708
rect 10534 -1714 10592 -1708
rect 10726 -1714 10784 -1708
rect 10918 -1714 10976 -1708
rect 11108 -1714 11166 -1708
rect 11304 -1716 11362 -1708
rect 11496 -1716 11554 -1708
rect 11688 -1712 11746 -1708
rect 6680 -1718 8458 -1716
rect 6680 -1726 6732 -1718
rect 6872 -1724 6924 -1718
rect 7064 -1724 7116 -1718
rect 7256 -1724 7308 -1718
rect 7448 -1724 7500 -1718
rect 7642 -1724 7694 -1718
rect 7832 -1724 7884 -1718
rect 8022 -1726 8074 -1718
rect 8212 -1722 8270 -1718
rect 8406 -1722 8458 -1718
rect 5086 -2164 5226 -2050
rect 5022 -2166 5226 -2164
rect 5278 -2164 5418 -2050
rect 5606 -2050 5658 -2040
rect 5800 -2050 5954 -2040
rect 5992 -2050 6044 -2040
rect 6584 -2050 6636 -2040
rect 5470 -2164 5606 -2050
rect 5278 -2166 5606 -2164
rect 5658 -2166 5800 -2050
rect 5852 -2166 5992 -2050
rect 6044 -2166 6046 -2050
rect 6560 -2166 6584 -2056
rect 6776 -2050 6828 -2040
rect 6636 -2166 6776 -2056
rect 6970 -2050 7022 -2040
rect 6828 -2166 6970 -2056
rect 7162 -2052 7214 -2042
rect 7022 -2166 7162 -2056
rect 5034 -2174 5086 -2166
rect 5226 -2176 5278 -2166
rect 5418 -2174 5470 -2166
rect 5606 -2176 5658 -2166
rect 5800 -2176 5852 -2166
rect 5992 -2176 6044 -2166
rect 6584 -2176 6636 -2166
rect 6776 -2176 6828 -2166
rect 6970 -2176 7022 -2166
rect 7354 -2050 7406 -2040
rect 7214 -2166 7354 -2056
rect 7546 -2050 7598 -2040
rect 7406 -2166 7546 -2056
rect 7736 -2052 7788 -2042
rect 7598 -2166 7736 -2056
rect 7162 -2178 7214 -2168
rect 7354 -2176 7406 -2166
rect 7546 -2176 7598 -2166
rect 7928 -2050 7980 -2040
rect 7788 -2166 7928 -2056
rect 8120 -2050 8172 -2040
rect 7980 -2166 8120 -2056
rect 8212 -2056 8266 -1722
rect 9100 -2034 9152 -2030
rect 9288 -2034 9340 -2032
rect 9484 -2034 9536 -2032
rect 9674 -2034 9726 -2030
rect 9868 -2034 9920 -2030
rect 10058 -2034 10110 -2032
rect 10248 -2034 10300 -2032
rect 10442 -2034 10494 -2030
rect 10632 -2034 10684 -2032
rect 10826 -2034 10878 -2030
rect 11020 -2034 11072 -2030
rect 11210 -2034 11262 -2030
rect 11404 -2034 11456 -2030
rect 11592 -2034 11644 -2032
rect 11786 -2034 11838 -2032
rect 11876 -2034 11940 -1708
rect 11978 -2034 12030 -2028
rect 9090 -2038 12030 -2034
rect 9090 -2040 11978 -2038
rect 8312 -2050 8364 -2040
rect 8172 -2166 8312 -2056
rect 8506 -2050 8558 -2040
rect 8364 -2166 8506 -2056
rect 8558 -2166 8564 -2056
rect 9090 -2156 9100 -2040
rect 9152 -2042 9674 -2040
rect 9152 -2156 9288 -2042
rect 9090 -2158 9288 -2156
rect 9340 -2158 9484 -2042
rect 9536 -2156 9674 -2042
rect 9726 -2156 9868 -2040
rect 9920 -2042 10442 -2040
rect 9920 -2156 10058 -2042
rect 9536 -2158 10058 -2156
rect 10110 -2158 10248 -2042
rect 10300 -2156 10442 -2042
rect 10494 -2042 10826 -2040
rect 10494 -2156 10632 -2042
rect 10300 -2158 10632 -2156
rect 10684 -2156 10826 -2042
rect 10878 -2156 11020 -2040
rect 11072 -2156 11210 -2040
rect 11262 -2156 11404 -2040
rect 11456 -2042 11978 -2040
rect 11456 -2156 11592 -2042
rect 10684 -2158 11592 -2156
rect 11644 -2158 11786 -2042
rect 11838 -2154 11978 -2042
rect 11838 -2158 12030 -2154
rect 9090 -2162 12030 -2158
rect 9100 -2166 9152 -2162
rect 7736 -2178 7788 -2168
rect 7928 -2176 7980 -2166
rect 8120 -2176 8172 -2166
rect 8312 -2176 8364 -2166
rect 8506 -2176 8558 -2166
rect 9288 -2168 9340 -2162
rect 9484 -2168 9536 -2162
rect 9674 -2166 9726 -2162
rect 9868 -2166 9920 -2162
rect 10058 -2168 10110 -2162
rect 10248 -2168 10300 -2162
rect 10442 -2166 10494 -2162
rect 10632 -2168 10684 -2162
rect 10826 -2166 10878 -2162
rect 11020 -2166 11072 -2162
rect 11210 -2166 11262 -2162
rect 11404 -2166 11456 -2162
rect 11592 -2168 11644 -2162
rect 11786 -2168 11838 -2162
rect 11978 -2164 12030 -2162
rect 9194 -2498 9246 -2492
rect 9386 -2498 9438 -2492
rect 9578 -2498 9630 -2494
rect 9772 -2498 9824 -2492
rect 9960 -2498 10012 -2494
rect 10154 -2498 10206 -2494
rect 10344 -2498 10396 -2494
rect 10538 -2498 10590 -2494
rect 10730 -2498 10782 -2494
rect 10924 -2498 10976 -2492
rect 11112 -2498 11164 -2494
rect 11306 -2498 11358 -2492
rect 11498 -2498 11550 -2494
rect 11688 -2498 11740 -2492
rect 11884 -2498 11936 -2494
rect 4226 -2510 4278 -2500
rect 4416 -2510 4468 -2500
rect 4608 -2510 4660 -2502
rect 5128 -2506 5180 -2500
rect 5320 -2506 5372 -2500
rect 5514 -2506 5566 -2502
rect 5702 -2506 5754 -2500
rect 5898 -2506 5950 -2500
rect 5126 -2510 5950 -2506
rect 6680 -2510 6732 -2502
rect 6874 -2510 6926 -2502
rect 7066 -2510 7118 -2502
rect 7256 -2510 7308 -2502
rect 7448 -2510 7500 -2502
rect 7640 -2510 7692 -2504
rect 7834 -2510 7886 -2502
rect 8024 -2510 8076 -2502
rect 8216 -2510 8268 -2500
rect 9186 -2502 11940 -2498
rect 8408 -2510 8460 -2504
rect 4214 -2626 4226 -2510
rect 4278 -2626 4416 -2510
rect 4468 -2512 4670 -2510
rect 4468 -2626 4608 -2512
rect 4214 -2628 4608 -2626
rect 4660 -2628 4670 -2512
rect 5126 -2626 5128 -2510
rect 5180 -2626 5320 -2510
rect 5372 -2512 5702 -2510
rect 5372 -2626 5514 -2512
rect 5126 -2628 5514 -2626
rect 5566 -2626 5702 -2512
rect 5754 -2626 5898 -2510
rect 6672 -2512 8216 -2510
rect 6094 -2566 6164 -2556
rect 5950 -2620 6094 -2566
rect 5950 -2626 6164 -2620
rect 5566 -2628 5950 -2626
rect 4226 -2636 4278 -2628
rect 4416 -2636 4468 -2628
rect 4608 -2638 4660 -2628
rect 5128 -2636 5180 -2628
rect 5320 -2636 5372 -2628
rect 5514 -2638 5566 -2628
rect 5702 -2636 5754 -2628
rect 5898 -2636 5950 -2628
rect 6094 -2630 6164 -2626
rect 6672 -2628 6680 -2512
rect 6732 -2628 6874 -2512
rect 6926 -2628 7066 -2512
rect 7118 -2628 7256 -2512
rect 7308 -2628 7448 -2512
rect 7500 -2514 7834 -2512
rect 7500 -2628 7640 -2514
rect 6680 -2638 6732 -2628
rect 6874 -2638 6926 -2628
rect 7066 -2638 7118 -2628
rect 7256 -2638 7308 -2628
rect 7448 -2638 7500 -2628
rect 7692 -2628 7834 -2514
rect 7886 -2628 8024 -2512
rect 8076 -2626 8216 -2512
rect 8268 -2514 8464 -2510
rect 8268 -2626 8408 -2514
rect 8076 -2628 8408 -2626
rect 7640 -2640 7692 -2630
rect 7834 -2638 7886 -2628
rect 8024 -2638 8076 -2628
rect 8216 -2636 8268 -2628
rect 8460 -2572 8464 -2514
rect 8614 -2572 8678 -2562
rect 8460 -2626 8614 -2572
rect 9186 -2618 9194 -2502
rect 9246 -2618 9386 -2502
rect 9438 -2504 9772 -2502
rect 9438 -2618 9578 -2504
rect 9186 -2620 9578 -2618
rect 9630 -2618 9772 -2504
rect 9824 -2504 10924 -2502
rect 9824 -2618 9960 -2504
rect 9630 -2620 9960 -2618
rect 10012 -2620 10154 -2504
rect 10206 -2620 10344 -2504
rect 10396 -2620 10538 -2504
rect 10590 -2620 10730 -2504
rect 10782 -2618 10924 -2504
rect 10976 -2504 11306 -2502
rect 10976 -2618 11112 -2504
rect 10782 -2620 11112 -2618
rect 11164 -2618 11306 -2504
rect 11358 -2504 11688 -2502
rect 11358 -2618 11498 -2504
rect 11164 -2620 11498 -2618
rect 11550 -2618 11688 -2504
rect 11740 -2504 11940 -2502
rect 11740 -2618 11884 -2504
rect 11550 -2620 11884 -2618
rect 11936 -2556 11940 -2504
rect 12092 -2556 12148 -2548
rect 11936 -2558 12148 -2556
rect 11936 -2614 12092 -2558
rect 11936 -2620 11940 -2614
rect 9186 -2622 11940 -2620
rect 8460 -2628 8678 -2626
rect 9194 -2628 9246 -2622
rect 9386 -2628 9438 -2622
rect 8408 -2640 8460 -2630
rect 8614 -2636 8678 -2628
rect 9578 -2630 9630 -2622
rect 9772 -2628 9824 -2622
rect 9960 -2630 10012 -2622
rect 10154 -2630 10206 -2622
rect 10344 -2630 10396 -2622
rect 10538 -2630 10590 -2622
rect 10730 -2630 10782 -2622
rect 10924 -2628 10976 -2622
rect 11112 -2630 11164 -2622
rect 11306 -2628 11358 -2622
rect 11498 -2630 11550 -2622
rect 11688 -2628 11740 -2622
rect 11884 -2630 11936 -2622
rect 12092 -2624 12148 -2614
use sky130_fd_pr__nfet_01v8_42S873  XM1
timestamp 1709130382
transform 1 0 4491 0 1 -2038
box -407 -810 407 810
use sky130_fd_pr__pfet_01v8_UYM7GH  XM2
timestamp 1709130382
transform 1 0 4207 0 1 863
box -407 -2019 407 2019
use sky130_fd_pr__pfet_01v8_VC5S4W  XM3
timestamp 1709130382
transform 1 0 5807 0 1 2493
box -647 -1019 647 1019
use sky130_fd_pr__pfet_01v8_VC5S4W  XM4
timestamp 1709130382
transform 1 0 5541 0 1 189
box -647 -1019 647 1019
use sky130_fd_pr__nfet_01v8_JT8PYA  XM5
timestamp 1709130382
transform 1 0 5539 0 1 -2338
box -647 -510 647 510
use sky130_fd_pr__nfet_01v8_JLF2PR  XM6
timestamp 1709130382
transform -1 0 5539 0 1 -1424
box -647 -510 647 510
use sky130_fd_pr__pfet_01v8_VC5YSW  XM7
timestamp 1709130382
transform 1 0 7475 0 1 2493
box -1127 -1019 1127 1019
use sky130_fd_pr__pfet_01v8_VC5YSW  XM8
timestamp 1709130382
transform 1 0 7571 0 1 191
box -1127 -1019 1127 1019
use sky130_fd_pr__nfet_01v8_Z85QYA  XM9
timestamp 1709130382
transform 1 0 7571 0 1 -2340
box -1127 -510 1127 510
use sky130_fd_pr__nfet_01v8_PPAFLS  XM10
timestamp 1709130382
transform -1 0 7571 0 1 -1426
box -1127 -510 1127 510
use sky130_fd_pr__pfet_01v8_VC56GX  XM11
timestamp 1709130382
transform 1 0 10103 0 1 2493
box -1607 -1019 1607 1019
use sky130_fd_pr__pfet_01v8_VC56GX  XM12
timestamp 1709130382
transform 1 0 10565 0 1 191
box -1607 -1019 1607 1019
use sky130_fd_pr__nfet_01v8_CDSMYA  XM13
timestamp 1709130382
transform 1 0 10565 0 1 -2330
box -1607 -510 1607 510
use sky130_fd_pr__nfet_01v8_UBPJLS  XM14
timestamp 1709130382
transform -1 0 10565 0 1 -1416
box -1607 -510 1607 510
<< labels >>
flabel metal1 3796 -1476 3996 -1276 0 FreeSans 256 0 0 0 vctrl
port 2 nsew
flabel metal1 3828 -2844 4028 -2644 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal1 11970 -948 12170 -748 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 3798 3312 3998 3512 0 FreeSans 256 0 0 0 vdd
port 0 nsew
<< end >>
