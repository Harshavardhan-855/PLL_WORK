** sch_path: /home/harsh/design/xschem/PLL_FOLDER/cp/cp_schem.sch
.subckt cp_schem vdd cp_bias qa cp_out qb vss
*.PININFO qa:I qb:I cp_out:O vdd:B vss:B cp_bias:I
XM1 n1 n1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=6 nf=3 m=1
XM2 n1 bias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=2 nf=2 m=1
XM3 bias bias vss vss sky130_fd_pr__nfet_01v8 L=0.30 W=2 nf=2 m=1
XM4 n2 n1 vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=14 nf=7 m=1
XM5 n3 bias vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=0.7 nf=1 m=1
XM6 cp_out qa n2 vdd sky130_fd_pr__pfet_01v8 L=2 W=1 nf=1 m=1
XM7 cp_out qb n3 vss sky130_fd_pr__nfet_01v8 L=5 W=1 nf=1 m=1
XM8 bias cp_bias vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=18 nf=9 m=1
.ends
.end
